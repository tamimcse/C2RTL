`include "component_library.v"
`include "macros.v"

`timescale 1ns / 1ps
module top(clock, sb_subset_123_D, sbbit6_121_D, sbbit5_120_D, sbbit4_119_D, sbbit3_118_D, sbbit2_117_D, sbbit1_116_D, bs_subset_114_D, bsbit6_112_D, bsbit5_111_D, bsbit4_110_D, bsbit3_109_D, bsbit2_108_D, bsbit1_107_D, ss_subset_104_D, ssbit6_102_D, ssbit5_101_D, ssbit4_100_D, ip_dst_99_D, ssbit3_98_D, ssbit2_97_D, ssbit1_96_D, ip_src_95_D, R149);
  //IN
  input clock;
  input [63:0] sb_subset_123_D;
  input [31:0] sbbit6_121_D;
  input [31:0] sbbit5_120_D;
  input [31:0] sbbit4_119_D;
  input [31:0] sbbit3_118_D;
  input [31:0] sbbit2_117_D;
  input [31:0] sbbit1_116_D;
  input [63:0] bs_subset_114_D;
  input [31:0] bsbit6_112_D;
  input [31:0] bsbit5_111_D;
  input [31:0] bsbit4_110_D;
  input [31:0] bsbit3_109_D;
  input [31:0] bsbit2_108_D;
  input [31:0] bsbit1_107_D;
  input [63:0] ss_subset_104_D;
  input [31:0] ssbit6_102_D;
  input [31:0] ssbit5_101_D;
  input [31:0] ssbit4_100_D;
  input [31:0] ip_dst_99_D;
  input [31:0] ssbit3_98_D;
  input [31:0] ssbit2_97_D;
  input [31:0] ssbit1_96_D;
  input [31:0] ip_src_95_D;
  //OUT
  output [15:0] R149;
  //WIRES
  wire [15:0] R149;
  wire [31:0] R148;
  wire [31:0] R147;
  wire [31:0] R146;
  wire [63:0] R145;
  wire [63:0] R144;
  wire [63:0] R143;
  wire [63:0] R142;
  wire [63:0] R141;
  wire [63:0] R140;
  wire [15:0] R139;
  wire [15:0] R138;
  wire [15:0] R137;
  wire [15:0] R136;
  wire [15:0] R135;
  wire [15:0] R134;
  wire [15:0] R133;
  wire [15:0] R132;
  wire [15:0] R131;
  wire [15:0] R130;
  wire [15:0] R129;
  wire [15:0] R128;
  wire [15:0] R127;
  wire [15:0] R126;
  wire [15:0] R125;
  wire [31:0] R124;
  wire [31:0] R123;
  wire [31:0] R122;
  wire [31:0] R121;
  wire [31:0] R120;
  wire [31:0] R119;
  wire [31:0] R118;
  wire [31:0] R117;
  wire [31:0] R116;
  wire [15:0] mux2;
  wire [15:0] mux1;
  wire [15:0] mux0;
  wire [15:0] _131;
  wire [15:0] _132;
  wire [0:0] ifout109;
  wire [15:0] _133;
  wire [15:0] _134;
  wire [0:0] ifout106;
  wire [0:0] ifout105;
  wire [15:0] sb_matchid_130;
  wire [31:0] _93;
  wire [15:0] sb_priority_129;
  wire [15:0] bs_matchid_128;
  wire [31:0] _92;
  wire [15:0] bs_priority_127;
  wire [15:0] ss_matchid_126;
  wire [31:0] _91;
  wire [15:0] ss_priority_125;
  wire [31:0] sb_leaf_124;
  wire [63:0] _90;
  wire [63:0] _89;
  wire [63:0] _88;
  wire [15:0] sb_idx_122;
  wire [15:0] _87;
  wire [15:0] _86;
  wire [15:0] _85;
  wire [31:0] _84;
  wire [15:0] _83;
  wire [15:0] _82;
  wire [15:0] _81;
  wire [15:0] _80;
  wire [31:0] _79;
  wire [15:0] _78;
  wire [15:0] _77;
  wire [15:0] _76;
  wire [15:0] _75;
  wire [31:0] _74;
  wire [15:0] _73;
  wire [15:0] _72;
  wire [15:0] _71;
  wire [15:0] _70;
  wire [31:0] _69;
  wire [15:0] _68;
  wire [15:0] _67;
  wire [15:0] _66;
  wire [15:0] _65;
  wire [31:0] _64;
  wire [15:0] _63;
  wire [15:0] _62;
  wire [31:0] _61;
  wire [31:0] bs_leaf_115;
  wire [63:0] _60;
  wire [63:0] _59;
  wire [63:0] _58;
  wire [15:0] bs_idx_113;
  wire [15:0] _57;
  wire [15:0] _56;
  wire [15:0] _55;
  wire [31:0] _54;
  wire [15:0] _53;
  wire [15:0] _52;
  wire [15:0] _51;
  wire [15:0] _50;
  wire [31:0] _49;
  wire [15:0] _48;
  wire [15:0] _47;
  wire [15:0] _46;
  wire [15:0] _45;
  wire [31:0] _44;
  wire [15:0] _43;
  wire [15:0] _42;
  wire [15:0] _41;
  wire [15:0] _40;
  wire [31:0] _39;
  wire [15:0] _38;
  wire [15:0] _37;
  wire [15:0] _36;
  wire [15:0] _35;
  wire [31:0] _34;
  wire [15:0] _33;
  wire [15:0] _32;
  wire [31:0] _31;
  wire [31:0] ss_leaf_106;
  wire [63:0] _30;
  wire [63:0] _29;
  wire [63:0] _28;
  wire [15:0] ss_idx_103;
  wire [15:0] _27;
  wire [15:0] _26;
  wire [15:0] _25;
  wire [31:0] _24;
  wire [15:0] _23;
  wire [15:0] _22;
  wire [15:0] _21;
  wire [15:0] _20;
  wire [31:0] _19;
  wire [15:0] _18;
  wire [15:0] _17;
  wire [15:0] _16;
  wire [15:0] _15;
  wire [31:0] _14;
  wire [15:0] _13;
  wire [15:0] _12;
  wire [15:0] _11;
  wire [15:0] _10;
  wire [31:0] _9;
  wire [15:0] _8;
  wire [15:0] _7;
  wire [15:0] _6;
  wire [15:0] _5;
  wire [31:0] _4;
  wire [15:0] _3;
  wire [15:0] _2;
  wire [31:0] _1;
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op72 (.out1(_69), .in1(ip_src_95_D), .in2(sbbit3_118_D));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op67 (.out1(_64), .in1(ip_src_95_D), .in2(sbbit2_117_D));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op40 (.out1(_39), .in1(ip_dst_99_D), .in2(bsbit3_109_D));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op35 (.out1(_34), .in1(ip_dst_99_D), .in2(bsbit2_108_D));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op8 (.out1(_9), .in1(ip_src_95_D), .in2(ssbit3_98_D));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op3 (.out1(_4), .in1(ip_src_95_D), .in2(ssbit2_97_D));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op87 (.out1(_84), .in1(ip_src_95_D), .in2(sbbit6_121_D));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op82 (.out1(_79), .in1(ip_src_95_D), .in2(sbbit5_120_D));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op77 (.out1(_74), .in1(ip_src_95_D), .in2(sbbit4_119_D));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op55 (.out1(_54), .in1(ip_dst_99_D), .in2(bsbit6_112_D));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op50 (.out1(_49), .in1(ip_dst_99_D), .in2(bsbit5_111_D));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op45 (.out1(_44), .in1(ip_dst_99_D), .in2(bsbit4_110_D));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op23 (.out1(_24), .in1(ip_dst_99_D), .in2(ssbit6_102_D));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op18 (.out1(_19), .in1(ip_dst_99_D), .in2(ssbit5_101_D));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op13 (.out1(_14), .in1(ip_dst_99_D), .in2(ssbit4_100_D));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op73 (.out1(_70), .in1(_69));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op68 (.out1(_65), .in1(_64));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op41 (.out1(_40), .in1(_39));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op36 (.out1(_35), .in1(_34));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op9 (.out1(_10), .in1(_9));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op4 (.out1(_5), .in1(_4));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op115 (.out1(R116), .clock(clock), .in1(_84));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op116 (.out1(R117), .clock(clock), .in1(_79));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op117 (.out1(R118), .clock(clock), .in1(_74));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op118 (.out1(R119), .clock(clock), .in1(_54));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op119 (.out1(R120), .clock(clock), .in1(_49));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op120 (.out1(R121), .clock(clock), .in1(_44));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op121 (.out1(R122), .clock(clock), .in1(_24));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op122 (.out1(R123), .clock(clock), .in1(_19));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op123 (.out1(R124), .clock(clock), .in1(_14));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op124 (.out1(R125), .clock(clock), .in1(_70));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op125 (.out1(R126), .clock(clock), .in1(_65));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op126 (.out1(R127), .clock(clock), .in1(_40));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op127 (.out1(R128), .clock(clock), .in1(_35));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op128 (.out1(R129), .clock(clock), .in1(_10));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op129 (.out1(R130), .clock(clock), .in1(_5));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op78 (.out1(_75), .in1(R118));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op46 (.out1(_45), .in1(R121));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op14 (.out1(_15), .in1(R124));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op83 (.out1(_80), .in1(R117));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op51 (.out1(_50), .in1(R120));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op19 (.out1(_20), .in1(R123));
  LSHIFT_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(1), .BITSIZE_out1(16), .PRECISION(16)) op69 (.out1(_66), .in1(R126), .in2(1 'd 1));
  LSHIFT_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(1), .BITSIZE_out1(16), .PRECISION(16)) op37 (.out1(_36), .in1(R128), .in2(1 'd 1));
  LSHIFT_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(1), .BITSIZE_out1(16), .PRECISION(16)) op5 (.out1(_6), .in1(R130), .in2(1 'd 1));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op88 (.out1(_85), .in1(R116));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op56 (.out1(_55), .in1(R119));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op24 (.out1(_25), .in1(R122));
  LSHIFT_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(2), .BITSIZE_out1(16), .PRECISION(16)) op74 (.out1(_71), .in1(R125), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(2), .BITSIZE_out1(16), .PRECISION(16)) op42 (.out1(_41), .in1(R127), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(2), .BITSIZE_out1(16), .PRECISION(16)) op10 (.out1(_11), .in1(R129), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(2), .BITSIZE_out1(16), .PRECISION(16)) op79 (.out1(_76), .in1(_75), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(2), .BITSIZE_out1(16), .PRECISION(16)) op47 (.out1(_46), .in1(_45), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(2), .BITSIZE_out1(16), .PRECISION(16)) op15 (.out1(_16), .in1(_15), .in2(2 'd 3));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op64 (.out1(_61), .in1(ip_src_95_D), .in2(sbbit1_116_D));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op32 (.out1(_31), .in1(ip_dst_99_D), .in2(bsbit1_107_D));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op0 (.out1(_1), .in1(ip_src_95_D), .in2(ssbit1_96_D));
  LSHIFT_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(3), .BITSIZE_out1(16), .PRECISION(16)) op84 (.out1(_81), .in1(_80), .in2(3 'd 4));
  LSHIFT_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(3), .BITSIZE_out1(16), .PRECISION(16)) op52 (.out1(_51), .in1(_50), .in2(3 'd 4));
  LSHIFT_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(3), .BITSIZE_out1(16), .PRECISION(16)) op20 (.out1(_21), .in1(_20), .in2(3 'd 4));
  LSHIFT_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(3), .BITSIZE_out1(16), .PRECISION(16)) op89 (.out1(_86), .in1(_85), .in2(3 'd 5));
  LSHIFT_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(3), .BITSIZE_out1(16), .PRECISION(16)) op57 (.out1(_56), .in1(_55), .in2(3 'd 5));
  LSHIFT_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(3), .BITSIZE_out1(16), .PRECISION(16)) op25 (.out1(_26), .in1(_25), .in2(3 'd 5));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op65 (.out1(_62), .in1(_61));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op33 (.out1(_32), .in1(_31));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op1 (.out1(_2), .in1(_1));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(2), .BITSIZE_out1(16)) op70 (.out1(_67), .in1(_66), .in2(2 'd 2));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(1), .BITSIZE_out1(16)) op66 (.out1(_63), .in1(_62), .in2(1 'd 1));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(2), .BITSIZE_out1(16)) op38 (.out1(_37), .in1(_36), .in2(2 'd 2));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(1), .BITSIZE_out1(16)) op34 (.out1(_33), .in1(_32), .in2(1 'd 1));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(2), .BITSIZE_out1(16)) op6 (.out1(_7), .in1(_6), .in2(2 'd 2));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(1), .BITSIZE_out1(16)) op2 (.out1(_3), .in1(_2), .in2(1 'd 1));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(3), .BITSIZE_out1(16)) op75 (.out1(_72), .in1(_71), .in2(3 'd 4));
  bit_or #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op71 (.out1(_68), .in1(_63), .in2(_67));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(3), .BITSIZE_out1(16)) op43 (.out1(_42), .in1(_41), .in2(3 'd 4));
  bit_or #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op39 (.out1(_38), .in1(_33), .in2(_37));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(3), .BITSIZE_out1(16)) op11 (.out1(_12), .in1(_11), .in2(3 'd 4));
  bit_or #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op7 (.out1(_8), .in1(_3), .in2(_7));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(4), .BITSIZE_out1(16)) op80 (.out1(_77), .in1(_76), .in2(4 'd 8));
  bit_or #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op76 (.out1(_73), .in1(_68), .in2(_72));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(4), .BITSIZE_out1(16)) op48 (.out1(_47), .in1(_46), .in2(4 'd 8));
  bit_or #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op44 (.out1(_43), .in1(_38), .in2(_42));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(4), .BITSIZE_out1(16)) op16 (.out1(_17), .in1(_16), .in2(4 'd 8));
  bit_or #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op12 (.out1(_13), .in1(_8), .in2(_12));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(5), .BITSIZE_out1(16)) op85 (.out1(_82), .in1(_81), .in2(5 'd 16));
  bit_or #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op81 (.out1(_78), .in1(_73), .in2(_77));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(5), .BITSIZE_out1(16)) op53 (.out1(_52), .in1(_51), .in2(5 'd 16));
  bit_or #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op49 (.out1(_48), .in1(_43), .in2(_47));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(5), .BITSIZE_out1(16)) op21 (.out1(_22), .in1(_21), .in2(5 'd 16));
  bit_or #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op17 (.out1(_18), .in1(_13), .in2(_17));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op130 (.out1(R131), .clock(clock), .in1(_86));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op131 (.out1(R132), .clock(clock), .in1(_56));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op132 (.out1(R133), .clock(clock), .in1(_26));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op133 (.out1(R134), .clock(clock), .in1(_82));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op134 (.out1(R135), .clock(clock), .in1(_78));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op135 (.out1(R136), .clock(clock), .in1(_52));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op136 (.out1(R137), .clock(clock), .in1(_48));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op137 (.out1(R138), .clock(clock), .in1(_22));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op138 (.out1(R139), .clock(clock), .in1(_18));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(6), .BITSIZE_out1(16)) op90 (.out1(_87), .in1(R131), .in2(6 'd 32));
  bit_or #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op86 (.out1(_83), .in1(R135), .in2(R134));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(6), .BITSIZE_out1(16)) op58 (.out1(_57), .in1(R132), .in2(6 'd 32));
  bit_or #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op54 (.out1(_53), .in1(R137), .in2(R136));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(6), .BITSIZE_out1(16)) op26 (.out1(_27), .in1(R133), .in2(6 'd 32));
  bit_or #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op22 (.out1(_23), .in1(R139), .in2(R138));
  bit_or #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op91 (.out1(sb_idx_122), .in1(_83), .in2(_87));
  bit_or #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op59 (.out1(bs_idx_113), .in1(_53), .in2(_57));
  bit_or #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op27 (.out1(ss_idx_103), .in1(_23), .in2(_27));
  cast #(.BITSIZE_in1(16), .BITSIZE_out1(64)) op92 (.out1(_88), .in1(sb_idx_122));
  cast #(.BITSIZE_in1(16), .BITSIZE_out1(64)) op60 (.out1(_58), .in1(bs_idx_113));
  cast #(.BITSIZE_in1(16), .BITSIZE_out1(64)) op28 (.out1(_28), .in1(ss_idx_103));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op93 (.out1(_89), .in1(_88), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op61 (.out1(_59), .in1(_58), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op29 (.out1(_29), .in1(_28), .in2(2 'd 2));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op139 (.out1(R140), .clock(clock), .in1(_89));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op140 (.out1(R141), .clock(clock), .in1(_59));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op141 (.out1(R142), .clock(clock), .in1(_29));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op94 (.out1(_90), .in1(sb_subset_123_D), .in2(R140));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op62 (.out1(_60), .in1(bs_subset_114_D), .in2(R141));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op30 (.out1(_30), .in1(ss_subset_104_D), .in2(R142));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op142 (.out1(R143), .clock(clock), .in1(_90));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op143 (.out1(R144), .clock(clock), .in1(_60));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op144 (.out1(R145), .clock(clock), .in1(_30));
  SRAM op95 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(sb_leaf_124),.ADR(R143));
  SRAM op63 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(bs_leaf_115),.ADR(R144));
  SRAM op31 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(ss_leaf_106),.ADR(R145));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op145 (.out1(R146), .clock(clock), .in1(sb_leaf_124));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op146 (.out1(R147), .clock(clock), .in1(bs_leaf_115));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op147 (.out1(R148), .clock(clock), .in1(ss_leaf_106));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(5), .BITSIZE_out1(32), .PRECISION(32)) op103 (.out1(_93), .in1(R146), .in2(5 'd 16));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(5), .BITSIZE_out1(32), .PRECISION(32)) op100 (.out1(_92), .in1(R147), .in2(5 'd 16));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(5), .BITSIZE_out1(32), .PRECISION(32)) op97 (.out1(_91), .in1(R148), .in2(5 'd 16));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op99 (.out1(bs_priority_127), .in1(R147));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op96 (.out1(ss_priority_125), .in1(R148));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op102 (.out1(sb_priority_129), .in1(R146));
  GT_EXPR #(.BITSIZE_in1(16), .BITSIZE_in2(16),.BITSIZE_out1(1)) op105 (.out1(ifout105), .in1(ss_priority_125), .in2(bs_priority_127));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op104 (.out1(sb_matchid_130), .in1(_93));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op101 (.out1(bs_matchid_128), .in1(_92));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op98 (.out1(ss_matchid_126), .in1(_91));
  GT_EXPR #(.BITSIZE_in1(16), .BITSIZE_in2(16),.BITSIZE_out1(1)) op109 (.out1(ifout109), .in1(bs_priority_127), .in2(sb_priority_129));
  GT_EXPR #(.BITSIZE_in1(16), .BITSIZE_in2(16),.BITSIZE_out1(1)) op106 (.out1(ifout106), .in1(ss_priority_125), .in2(sb_priority_129));
  assignment #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op111 (.out1(_131), .in1(sb_matchid_130));
  assignment #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op110 (.out1(_132), .in1(bs_matchid_128));
  assignment #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op108 (.out1(_133), .in1(sb_matchid_130));
  assignment #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op107 (.out1(_134), .in1(ss_matchid_126));
  MUX_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op112 (.out1(mux0), .in1(_131), .in2(_132), .sel(ifout109));
  MUX_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op113 (.out1(mux1), .in1(_133), .in2(_134), .sel(ifout106));
  MUX_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op114 (.out1(mux2), .in1(mux0), .in2(mux1), .sel(ifout105));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op148 (.out1(R149), .clock(clock), .in1(mux2));
endmodule