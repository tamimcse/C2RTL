`include "component_library.v"
`include "macros.v"

`timescale 1ns / 1ps
module top(clock, sb_subset_141_D, sbbit6_139_D, sbbit5_138_D, sbbit4_137_D, sbbit3_136_D, sbbit2_135_D, sbbit1_134_D, bs_subset_132_D, bsbit6_130_D, bsbit5_129_D, bsbit4_128_D, bsbit3_127_D, bsbit2_126_D, bsbit1_125_D, ss_subset_122_D, ssbit6_120_D, ssbit5_119_D, ip_dst_118_D, ssbit4_117_D, ssbit3_116_D, ssbit2_115_D, ip_src_114_D, ssbit1_113_D, R167);
  //IN
  input clock;
  input [63:0] sb_subset_141_D;
  input [7:0] sbbit6_139_D;
  input [7:0] sbbit5_138_D;
  input [7:0] sbbit4_137_D;
  input [7:0] sbbit3_136_D;
  input [7:0] sbbit2_135_D;
  input [7:0] sbbit1_134_D;
  input [63:0] bs_subset_132_D;
  input [7:0] bsbit6_130_D;
  input [7:0] bsbit5_129_D;
  input [7:0] bsbit4_128_D;
  input [7:0] bsbit3_127_D;
  input [7:0] bsbit2_126_D;
  input [7:0] bsbit1_125_D;
  input [63:0] ss_subset_122_D;
  input [7:0] ssbit6_120_D;
  input [7:0] ssbit5_119_D;
  input [31:0] ip_dst_118_D;
  input [7:0] ssbit4_117_D;
  input [7:0] ssbit3_116_D;
  input [7:0] ssbit2_115_D;
  input [31:0] ip_src_114_D;
  input [7:0] ssbit1_113_D;
  //OUT
  output [15:0] R167;
  //WIRES
  wire [15:0] R167;
  wire [31:0] R166;
  wire [31:0] R165;
  wire [31:0] R164;
  wire [63:0] R163;
  wire [63:0] R162;
  wire [63:0] R161;
  wire [63:0] R160;
  wire [63:0] R159;
  wire [63:0] R158;
  wire [15:0] R157;
  wire [15:0] R156;
  wire [15:0] R155;
  wire [15:0] R154;
  wire [15:0] R153;
  wire [15:0] R152;
  wire [15:0] R151;
  wire [15:0] R150;
  wire [15:0] R149;
  wire [15:0] R148;
  wire [15:0] R147;
  wire [15:0] R146;
  wire [15:0] R145;
  wire [15:0] R144;
  wire [15:0] R143;
  wire [31:0] R142;
  wire [31:0] R141;
  wire [31:0] R140;
  wire [31:0] R139;
  wire [31:0] R138;
  wire [31:0] R137;
  wire [31:0] R136;
  wire [31:0] R135;
  wire [31:0] R134;
  wire [15:0] mux2;
  wire [15:0] mux1;
  wire [15:0] mux0;
  wire [15:0] _149;
  wire [15:0] _150;
  wire [0:0] ifout127;
  wire [15:0] _151;
  wire [15:0] _152;
  wire [0:0] ifout124;
  wire [0:0] ifout123;
  wire [15:0] sb_matchid_148;
  wire [31:0] _111;
  wire [15:0] sb_priority_147;
  wire [15:0] bs_matchid_146;
  wire [31:0] _110;
  wire [15:0] bs_priority_145;
  wire [15:0] ss_matchid_144;
  wire [31:0] _109;
  wire [15:0] ss_priority_143;
  wire [31:0] sb_leaf_142;
  wire [63:0] _108;
  wire [63:0] _107;
  wire [63:0] _106;
  wire [15:0] sb_idx_140;
  wire [15:0] _105;
  wire [15:0] _104;
  wire [15:0] _103;
  wire [31:0] _102;
  wire [31:0] _101;
  wire [15:0] _100;
  wire [15:0] _99;
  wire [15:0] _98;
  wire [15:0] _97;
  wire [31:0] _96;
  wire [31:0] _95;
  wire [15:0] _94;
  wire [15:0] _93;
  wire [15:0] _92;
  wire [15:0] _91;
  wire [31:0] _90;
  wire [31:0] _89;
  wire [15:0] _88;
  wire [15:0] _87;
  wire [15:0] _86;
  wire [15:0] _85;
  wire [31:0] _84;
  wire [31:0] _83;
  wire [15:0] _82;
  wire [15:0] _81;
  wire [15:0] _80;
  wire [15:0] _79;
  wire [31:0] _78;
  wire [31:0] _77;
  wire [15:0] _76;
  wire [15:0] _75;
  wire [31:0] _74;
  wire [31:0] _73;
  wire [31:0] bs_leaf_133;
  wire [63:0] _72;
  wire [63:0] _71;
  wire [63:0] _70;
  wire [15:0] bs_idx_131;
  wire [15:0] _69;
  wire [15:0] _68;
  wire [15:0] _67;
  wire [31:0] _66;
  wire [31:0] _65;
  wire [15:0] _64;
  wire [15:0] _63;
  wire [15:0] _62;
  wire [15:0] _61;
  wire [31:0] _60;
  wire [31:0] _59;
  wire [15:0] _58;
  wire [15:0] _57;
  wire [15:0] _56;
  wire [15:0] _55;
  wire [31:0] _54;
  wire [31:0] _53;
  wire [15:0] _52;
  wire [15:0] _51;
  wire [15:0] _50;
  wire [15:0] _49;
  wire [31:0] _48;
  wire [31:0] _47;
  wire [15:0] _46;
  wire [15:0] _45;
  wire [15:0] _44;
  wire [15:0] _43;
  wire [31:0] _42;
  wire [31:0] _41;
  wire [15:0] _40;
  wire [15:0] _39;
  wire [31:0] _38;
  wire [31:0] _37;
  wire [31:0] ss_leaf_124;
  wire [63:0] _36;
  wire [63:0] _35;
  wire [63:0] _34;
  wire [15:0] ss_idx_121;
  wire [15:0] _33;
  wire [15:0] _32;
  wire [15:0] _31;
  wire [31:0] _30;
  wire [31:0] _29;
  wire [15:0] _28;
  wire [15:0] _27;
  wire [15:0] _26;
  wire [15:0] _25;
  wire [31:0] _24;
  wire [31:0] _23;
  wire [15:0] _22;
  wire [15:0] _21;
  wire [15:0] _20;
  wire [15:0] _19;
  wire [31:0] _18;
  wire [31:0] _17;
  wire [15:0] _16;
  wire [15:0] _15;
  wire [15:0] _14;
  wire [15:0] _13;
  wire [31:0] _12;
  wire [31:0] _11;
  wire [15:0] _10;
  wire [15:0] _9;
  wire [15:0] _8;
  wire [15:0] _7;
  wire [31:0] _6;
  wire [31:0] _5;
  wire [15:0] _4;
  wire [15:0] _3;
  wire [31:0] _2;
  wire [31:0] _1;
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(32)) op86 (.out1(_83), .in1(sbbit3_136_D));
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(32)) op80 (.out1(_77), .in1(sbbit2_135_D));
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(32)) op48 (.out1(_47), .in1(bsbit3_127_D));
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(32)) op42 (.out1(_41), .in1(bsbit2_126_D));
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(32)) op10 (.out1(_11), .in1(ssbit3_116_D));
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(32)) op4 (.out1(_5), .in1(ssbit2_115_D));
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(32)) op104 (.out1(_101), .in1(sbbit6_139_D));
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(32)) op98 (.out1(_95), .in1(sbbit5_138_D));
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(32)) op92 (.out1(_89), .in1(sbbit4_137_D));
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(32)) op66 (.out1(_65), .in1(bsbit6_130_D));
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(32)) op60 (.out1(_59), .in1(bsbit5_129_D));
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(32)) op54 (.out1(_53), .in1(bsbit4_128_D));
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(32)) op28 (.out1(_29), .in1(ssbit6_120_D));
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(32)) op22 (.out1(_23), .in1(ssbit5_119_D));
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(32)) op16 (.out1(_17), .in1(ssbit4_117_D));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op87 (.out1(_84), .in1(ip_src_114_D), .in2(_83));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op81 (.out1(_78), .in1(ip_src_114_D), .in2(_77));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op49 (.out1(_48), .in1(ip_dst_118_D), .in2(_47));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op43 (.out1(_42), .in1(ip_dst_118_D), .in2(_41));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op11 (.out1(_12), .in1(ip_src_114_D), .in2(_11));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op5 (.out1(_6), .in1(ip_src_114_D), .in2(_5));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op105 (.out1(_102), .in1(ip_src_114_D), .in2(_101));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op99 (.out1(_96), .in1(ip_src_114_D), .in2(_95));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op93 (.out1(_90), .in1(ip_src_114_D), .in2(_89));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op67 (.out1(_66), .in1(ip_dst_118_D), .in2(_65));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op61 (.out1(_60), .in1(ip_dst_118_D), .in2(_59));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op55 (.out1(_54), .in1(ip_dst_118_D), .in2(_53));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op29 (.out1(_30), .in1(ip_dst_118_D), .in2(_29));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op23 (.out1(_24), .in1(ip_dst_118_D), .in2(_23));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op17 (.out1(_18), .in1(ip_dst_118_D), .in2(_17));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op88 (.out1(_85), .in1(_84));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op82 (.out1(_79), .in1(_78));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op50 (.out1(_49), .in1(_48));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op44 (.out1(_43), .in1(_42));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op12 (.out1(_13), .in1(_12));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op6 (.out1(_7), .in1(_6));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op133 (.out1(R134), .clock(clock), .in1(_102));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op134 (.out1(R135), .clock(clock), .in1(_96));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op135 (.out1(R136), .clock(clock), .in1(_90));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op136 (.out1(R137), .clock(clock), .in1(_66));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op137 (.out1(R138), .clock(clock), .in1(_60));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op138 (.out1(R139), .clock(clock), .in1(_54));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op139 (.out1(R140), .clock(clock), .in1(_30));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op140 (.out1(R141), .clock(clock), .in1(_24));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op141 (.out1(R142), .clock(clock), .in1(_18));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op142 (.out1(R143), .clock(clock), .in1(_85));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op143 (.out1(R144), .clock(clock), .in1(_79));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op144 (.out1(R145), .clock(clock), .in1(_49));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op145 (.out1(R146), .clock(clock), .in1(_43));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op146 (.out1(R147), .clock(clock), .in1(_13));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op147 (.out1(R148), .clock(clock), .in1(_7));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op94 (.out1(_91), .in1(R136));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op56 (.out1(_55), .in1(R139));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op18 (.out1(_19), .in1(R142));
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(32)) op76 (.out1(_73), .in1(sbbit1_134_D));
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(32)) op38 (.out1(_37), .in1(bsbit1_125_D));
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(32)) op0 (.out1(_1), .in1(ssbit1_113_D));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op100 (.out1(_97), .in1(R135));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op62 (.out1(_61), .in1(R138));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op24 (.out1(_25), .in1(R141));
  LSHIFT_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(1), .BITSIZE_out1(16), .PRECISION(16)) op83 (.out1(_80), .in1(R144), .in2(1 'd 1));
  LSHIFT_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(1), .BITSIZE_out1(16), .PRECISION(16)) op45 (.out1(_44), .in1(R146), .in2(1 'd 1));
  LSHIFT_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(1), .BITSIZE_out1(16), .PRECISION(16)) op7 (.out1(_8), .in1(R148), .in2(1 'd 1));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op106 (.out1(_103), .in1(R134));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op68 (.out1(_67), .in1(R137));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op30 (.out1(_31), .in1(R140));
  LSHIFT_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(2), .BITSIZE_out1(16), .PRECISION(16)) op89 (.out1(_86), .in1(R143), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(2), .BITSIZE_out1(16), .PRECISION(16)) op51 (.out1(_50), .in1(R145), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(2), .BITSIZE_out1(16), .PRECISION(16)) op13 (.out1(_14), .in1(R147), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(2), .BITSIZE_out1(16), .PRECISION(16)) op95 (.out1(_92), .in1(_91), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(2), .BITSIZE_out1(16), .PRECISION(16)) op57 (.out1(_56), .in1(_55), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(2), .BITSIZE_out1(16), .PRECISION(16)) op19 (.out1(_20), .in1(_19), .in2(2 'd 3));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op77 (.out1(_74), .in1(ip_src_114_D), .in2(_73));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op39 (.out1(_38), .in1(ip_dst_118_D), .in2(_37));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op1 (.out1(_2), .in1(ip_src_114_D), .in2(_1));
  LSHIFT_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(3), .BITSIZE_out1(16), .PRECISION(16)) op101 (.out1(_98), .in1(_97), .in2(3 'd 4));
  LSHIFT_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(3), .BITSIZE_out1(16), .PRECISION(16)) op63 (.out1(_62), .in1(_61), .in2(3 'd 4));
  LSHIFT_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(3), .BITSIZE_out1(16), .PRECISION(16)) op25 (.out1(_26), .in1(_25), .in2(3 'd 4));
  LSHIFT_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(3), .BITSIZE_out1(16), .PRECISION(16)) op107 (.out1(_104), .in1(_103), .in2(3 'd 5));
  LSHIFT_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(3), .BITSIZE_out1(16), .PRECISION(16)) op69 (.out1(_68), .in1(_67), .in2(3 'd 5));
  LSHIFT_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(3), .BITSIZE_out1(16), .PRECISION(16)) op31 (.out1(_32), .in1(_31), .in2(3 'd 5));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op78 (.out1(_75), .in1(_74));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op40 (.out1(_39), .in1(_38));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op2 (.out1(_3), .in1(_2));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(2), .BITSIZE_out1(16)) op84 (.out1(_81), .in1(_80), .in2(2 'd 2));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(1), .BITSIZE_out1(16)) op79 (.out1(_76), .in1(_75), .in2(1 'd 1));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(2), .BITSIZE_out1(16)) op46 (.out1(_45), .in1(_44), .in2(2 'd 2));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(1), .BITSIZE_out1(16)) op41 (.out1(_40), .in1(_39), .in2(1 'd 1));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(2), .BITSIZE_out1(16)) op8 (.out1(_9), .in1(_8), .in2(2 'd 2));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(1), .BITSIZE_out1(16)) op3 (.out1(_4), .in1(_3), .in2(1 'd 1));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(3), .BITSIZE_out1(16)) op90 (.out1(_87), .in1(_86), .in2(3 'd 4));
  bit_or #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op85 (.out1(_82), .in1(_76), .in2(_81));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(3), .BITSIZE_out1(16)) op52 (.out1(_51), .in1(_50), .in2(3 'd 4));
  bit_or #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op47 (.out1(_46), .in1(_40), .in2(_45));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(3), .BITSIZE_out1(16)) op14 (.out1(_15), .in1(_14), .in2(3 'd 4));
  bit_or #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op9 (.out1(_10), .in1(_4), .in2(_9));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(4), .BITSIZE_out1(16)) op96 (.out1(_93), .in1(_92), .in2(4 'd 8));
  bit_or #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op91 (.out1(_88), .in1(_82), .in2(_87));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(4), .BITSIZE_out1(16)) op58 (.out1(_57), .in1(_56), .in2(4 'd 8));
  bit_or #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op53 (.out1(_52), .in1(_46), .in2(_51));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(4), .BITSIZE_out1(16)) op20 (.out1(_21), .in1(_20), .in2(4 'd 8));
  bit_or #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op15 (.out1(_16), .in1(_10), .in2(_15));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(5), .BITSIZE_out1(16)) op102 (.out1(_99), .in1(_98), .in2(5 'd 16));
  bit_or #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op97 (.out1(_94), .in1(_88), .in2(_93));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(5), .BITSIZE_out1(16)) op64 (.out1(_63), .in1(_62), .in2(5 'd 16));
  bit_or #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op59 (.out1(_58), .in1(_52), .in2(_57));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(5), .BITSIZE_out1(16)) op26 (.out1(_27), .in1(_26), .in2(5 'd 16));
  bit_or #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op21 (.out1(_22), .in1(_16), .in2(_21));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op148 (.out1(R149), .clock(clock), .in1(_104));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op149 (.out1(R150), .clock(clock), .in1(_68));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op150 (.out1(R151), .clock(clock), .in1(_32));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op151 (.out1(R152), .clock(clock), .in1(_99));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op152 (.out1(R153), .clock(clock), .in1(_94));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op153 (.out1(R154), .clock(clock), .in1(_63));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op154 (.out1(R155), .clock(clock), .in1(_58));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op155 (.out1(R156), .clock(clock), .in1(_27));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op156 (.out1(R157), .clock(clock), .in1(_22));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(6), .BITSIZE_out1(16)) op108 (.out1(_105), .in1(R149), .in2(6 'd 32));
  bit_or #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op103 (.out1(_100), .in1(R153), .in2(R152));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(6), .BITSIZE_out1(16)) op70 (.out1(_69), .in1(R150), .in2(6 'd 32));
  bit_or #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op65 (.out1(_64), .in1(R155), .in2(R154));
  bit_and #(.BITSIZE_in1(16), .BITSIZE_in2(6), .BITSIZE_out1(16)) op32 (.out1(_33), .in1(R151), .in2(6 'd 32));
  bit_or #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op27 (.out1(_28), .in1(R157), .in2(R156));
  bit_or #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op109 (.out1(sb_idx_140), .in1(_100), .in2(_105));
  bit_or #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op71 (.out1(bs_idx_131), .in1(_64), .in2(_69));
  bit_or #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op33 (.out1(ss_idx_121), .in1(_28), .in2(_33));
  cast #(.BITSIZE_in1(16), .BITSIZE_out1(64)) op110 (.out1(_106), .in1(sb_idx_140));
  cast #(.BITSIZE_in1(16), .BITSIZE_out1(64)) op72 (.out1(_70), .in1(bs_idx_131));
  cast #(.BITSIZE_in1(16), .BITSIZE_out1(64)) op34 (.out1(_34), .in1(ss_idx_121));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op111 (.out1(_107), .in1(_106), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op73 (.out1(_71), .in1(_70), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op35 (.out1(_35), .in1(_34), .in2(2 'd 2));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op157 (.out1(R158), .clock(clock), .in1(_107));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op158 (.out1(R159), .clock(clock), .in1(_71));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op159 (.out1(R160), .clock(clock), .in1(_35));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op112 (.out1(_108), .in1(sb_subset_141_D), .in2(R158));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op74 (.out1(_72), .in1(bs_subset_132_D), .in2(R159));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op36 (.out1(_36), .in1(ss_subset_122_D), .in2(R160));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op160 (.out1(R161), .clock(clock), .in1(_108));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op161 (.out1(R162), .clock(clock), .in1(_72));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op162 (.out1(R163), .clock(clock), .in1(_36));
  SRAM op113 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(sb_leaf_142),.ADR(R161));
  SRAM op75 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(bs_leaf_133),.ADR(R162));
  SRAM op37 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(ss_leaf_124),.ADR(R163));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op163 (.out1(R164), .clock(clock), .in1(sb_leaf_142));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op164 (.out1(R165), .clock(clock), .in1(bs_leaf_133));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op165 (.out1(R166), .clock(clock), .in1(ss_leaf_124));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(5), .BITSIZE_out1(32), .PRECISION(32)) op121 (.out1(_111), .in1(R164), .in2(5 'd 16));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(5), .BITSIZE_out1(32), .PRECISION(32)) op118 (.out1(_110), .in1(R165), .in2(5 'd 16));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(5), .BITSIZE_out1(32), .PRECISION(32)) op115 (.out1(_109), .in1(R166), .in2(5 'd 16));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op117 (.out1(bs_priority_145), .in1(R165));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op114 (.out1(ss_priority_143), .in1(R166));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op120 (.out1(sb_priority_147), .in1(R164));
  GT_EXPR #(.BITSIZE_in1(16), .BITSIZE_in2(16),.BITSIZE_out1(1)) op123 (.out1(ifout123), .in1(ss_priority_143), .in2(bs_priority_145));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op122 (.out1(sb_matchid_148), .in1(_111));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op119 (.out1(bs_matchid_146), .in1(_110));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op116 (.out1(ss_matchid_144), .in1(_109));
  GT_EXPR #(.BITSIZE_in1(16), .BITSIZE_in2(16),.BITSIZE_out1(1)) op127 (.out1(ifout127), .in1(bs_priority_145), .in2(sb_priority_147));
  GT_EXPR #(.BITSIZE_in1(16), .BITSIZE_in2(16),.BITSIZE_out1(1)) op124 (.out1(ifout124), .in1(ss_priority_143), .in2(sb_priority_147));
  assignment #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op129 (.out1(_149), .in1(sb_matchid_148));
  assignment #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op128 (.out1(_150), .in1(bs_matchid_146));
  assignment #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op126 (.out1(_151), .in1(sb_matchid_148));
  assignment #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op125 (.out1(_152), .in1(ss_matchid_144));
  MUX_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op130 (.out1(mux0), .in1(_149), .in2(_150), .sel(ifout127));
  MUX_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op131 (.out1(mux1), .in1(_151), .in2(_152), .sel(ifout124));
  MUX_GATE #(.BITSIZE_in1(16), .BITSIZE_in2(16), .BITSIZE_out1(16)) op132 (.out1(mux2), .in1(mux0), .in2(mux1), .sel(ifout123));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op166 (.out1(R167), .clock(clock), .in1(mux2));
endmodule