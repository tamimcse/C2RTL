`include "component_library.v"
`include "macros.v"

`timescale 1ns / 1ps
module top(clock, sb_subset_108_D, sbbit6_106_D, sbbit5_105_D, sbbit4_104_D, sbbit3_103_D, sbbit2_102_D, sbbit1_101_D, bs_subset_99_D, bsbit6_97_D, bsbit5_96_D, bsbit4_95_D, bsbit3_94_D, bsbit2_93_D, bsbit1_92_D, ss_subset_89_D, ssbit6_87_D, ssbit5_86_D, ssbit4_85_D, ip_dst_84_D, ssbit3_83_D, ssbit2_82_D, ssbit1_81_D, ip_src_80_D, R140);
  //IN
  input clock;
  input [63:0] sb_subset_108_D;
  input [31:0] sbbit6_106_D;
  input [31:0] sbbit5_105_D;
  input [31:0] sbbit4_104_D;
  input [31:0] sbbit3_103_D;
  input [31:0] sbbit2_102_D;
  input [31:0] sbbit1_101_D;
  input [63:0] bs_subset_99_D;
  input [31:0] bsbit6_97_D;
  input [31:0] bsbit5_96_D;
  input [31:0] bsbit4_95_D;
  input [31:0] bsbit3_94_D;
  input [31:0] bsbit2_93_D;
  input [31:0] bsbit1_92_D;
  input [63:0] ss_subset_89_D;
  input [31:0] ssbit6_87_D;
  input [31:0] ssbit5_86_D;
  input [31:0] ssbit4_85_D;
  input [31:0] ip_dst_84_D;
  input [31:0] ssbit3_83_D;
  input [31:0] ssbit2_82_D;
  input [31:0] ssbit1_81_D;
  input [31:0] ip_src_80_D;
  //OUT
  output [7:0] R140;
  //WIRES
  wire [7:0] R140;
  wire [31:0] R139;
  wire [31:0] R138;
  wire [31:0] R137;
  wire [63:0] R136;
  wire [63:0] R135;
  wire [63:0] R134;
  wire [63:0] R133;
  wire [63:0] R132;
  wire [63:0] R131;
  wire [31:0] R130;
  wire [31:0] R129;
  wire [31:0] R128;
  wire [31:0] R127;
  wire [31:0] R126;
  wire [31:0] R125;
  wire [31:0] R124;
  wire [31:0] R123;
  wire [31:0] R122;
  wire [31:0] R121;
  wire [31:0] R120;
  wire [31:0] R119;
  wire [31:0] R118;
  wire [31:0] R117;
  wire [31:0] R116;
  wire [31:0] R115;
  wire [31:0] R114;
  wire [31:0] R113;
  wire [31:0] R112;
  wire [31:0] R111;
  wire [31:0] R110;
  wire [31:0] R109;
  wire [31:0] R108;
  wire [31:0] R107;
  wire [31:0] R106;
  wire [31:0] R105;
  wire [31:0] R104;
  wire [31:0] R103;
  wire [31:0] R102;
  wire [31:0] R101;
  wire [7:0] mux2;
  wire [7:0] mux1;
  wire [7:0] mux0;
  wire [7:0] _116;
  wire [7:0] _117;
  wire [0:0] ifout94;
  wire [7:0] _118;
  wire [7:0] _119;
  wire [0:0] ifout91;
  wire [0:0] ifout90;
  wire [15:0] sb_matchid_115;
  wire [31:0] _78;
  wire [15:0] sb_priority_114;
  wire [15:0] bs_matchid_113;
  wire [31:0] _77;
  wire [15:0] bs_priority_112;
  wire [15:0] ss_matchid_111;
  wire [31:0] _76;
  wire [15:0] ss_priority_110;
  wire [31:0] sb_leaf_109;
  wire [63:0] _75;
  wire [63:0] _74;
  wire [63:0] _73;
  wire [31:0] sb_idx_107;
  wire [31:0] _72;
  wire [31:0] _71;
  wire [31:0] _70;
  wire [31:0] _69;
  wire [31:0] _68;
  wire [31:0] _67;
  wire [31:0] _66;
  wire [31:0] _65;
  wire [31:0] _64;
  wire [31:0] _63;
  wire [31:0] _62;
  wire [31:0] _61;
  wire [31:0] _60;
  wire [31:0] _59;
  wire [31:0] _58;
  wire [31:0] _57;
  wire [31:0] _56;
  wire [31:0] _55;
  wire [31:0] _54;
  wire [31:0] _53;
  wire [31:0] _52;
  wire [31:0] _51;
  wire [31:0] bs_leaf_100;
  wire [63:0] _50;
  wire [63:0] _49;
  wire [63:0] _48;
  wire [31:0] bs_idx_98;
  wire [31:0] _47;
  wire [31:0] _46;
  wire [31:0] _45;
  wire [31:0] _44;
  wire [31:0] _43;
  wire [31:0] _42;
  wire [31:0] _41;
  wire [31:0] _40;
  wire [31:0] _39;
  wire [31:0] _38;
  wire [31:0] _37;
  wire [31:0] _36;
  wire [31:0] _35;
  wire [31:0] _34;
  wire [31:0] _33;
  wire [31:0] _32;
  wire [31:0] _31;
  wire [31:0] _30;
  wire [31:0] _29;
  wire [31:0] _28;
  wire [31:0] _27;
  wire [31:0] _26;
  wire [31:0] ss_leaf_91;
  wire [63:0] _25;
  wire [63:0] _24;
  wire [63:0] _23;
  wire [31:0] ss_idx_88;
  wire [31:0] _22;
  wire [31:0] _21;
  wire [31:0] _20;
  wire [31:0] _19;
  wire [31:0] _18;
  wire [31:0] _17;
  wire [31:0] _16;
  wire [31:0] _15;
  wire [31:0] _14;
  wire [31:0] _13;
  wire [31:0] _12;
  wire [31:0] _11;
  wire [31:0] _10;
  wire [31:0] _9;
  wire [31:0] _8;
  wire [31:0] _7;
  wire [31:0] _6;
  wire [31:0] _5;
  wire [31:0] _4;
  wire [31:0] _3;
  wire [31:0] _2;
  wire [31:0] _1;
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op68 (.out1(_65), .in1(ip_src_80_D), .in2(sbbit5_105_D));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op64 (.out1(_61), .in1(ip_src_80_D), .in2(sbbit4_104_D));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op60 (.out1(_57), .in1(ip_src_80_D), .in2(sbbit3_103_D));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op56 (.out1(_53), .in1(ip_src_80_D), .in2(sbbit2_102_D));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op41 (.out1(_40), .in1(ip_dst_84_D), .in2(bsbit5_96_D));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op37 (.out1(_36), .in1(ip_dst_84_D), .in2(bsbit4_95_D));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op33 (.out1(_32), .in1(ip_dst_84_D), .in2(bsbit3_94_D));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op29 (.out1(_28), .in1(ip_dst_84_D), .in2(bsbit2_93_D));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op14 (.out1(_15), .in1(ip_dst_84_D), .in2(ssbit5_86_D));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op10 (.out1(_11), .in1(ip_dst_84_D), .in2(ssbit4_85_D));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op6 (.out1(_7), .in1(ip_src_80_D), .in2(ssbit3_83_D));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op2 (.out1(_3), .in1(ip_src_80_D), .in2(ssbit2_82_D));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op100 (.out1(R101), .clock(clock), .in1(_65));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op101 (.out1(R102), .clock(clock), .in1(_61));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op102 (.out1(R103), .clock(clock), .in1(_57));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op103 (.out1(R104), .clock(clock), .in1(_53));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op104 (.out1(R105), .clock(clock), .in1(_40));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op105 (.out1(R106), .clock(clock), .in1(_36));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op106 (.out1(R107), .clock(clock), .in1(_32));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op107 (.out1(R108), .clock(clock), .in1(_28));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op108 (.out1(R109), .clock(clock), .in1(_15));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op109 (.out1(R110), .clock(clock), .in1(_11));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op110 (.out1(R111), .clock(clock), .in1(_7));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op111 (.out1(R112), .clock(clock), .in1(_3));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(3), .BITSIZE_out1(32), .PRECISION(32)) op69 (.out1(_66), .in1(R101), .in2(3 'd 4));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(2), .BITSIZE_out1(32), .PRECISION(32)) op65 (.out1(_62), .in1(R102), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(2), .BITSIZE_out1(32), .PRECISION(32)) op61 (.out1(_58), .in1(R103), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(1), .BITSIZE_out1(32), .PRECISION(32)) op57 (.out1(_54), .in1(R104), .in2(1 'd 1));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(3), .BITSIZE_out1(32), .PRECISION(32)) op42 (.out1(_41), .in1(R105), .in2(3 'd 4));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(2), .BITSIZE_out1(32), .PRECISION(32)) op38 (.out1(_37), .in1(R106), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(2), .BITSIZE_out1(32), .PRECISION(32)) op34 (.out1(_33), .in1(R107), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(1), .BITSIZE_out1(32), .PRECISION(32)) op30 (.out1(_29), .in1(R108), .in2(1 'd 1));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(3), .BITSIZE_out1(32), .PRECISION(32)) op15 (.out1(_16), .in1(R109), .in2(3 'd 4));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(2), .BITSIZE_out1(32), .PRECISION(32)) op11 (.out1(_12), .in1(R110), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(2), .BITSIZE_out1(32), .PRECISION(32)) op7 (.out1(_8), .in1(R111), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(1), .BITSIZE_out1(32), .PRECISION(32)) op3 (.out1(_4), .in1(R112), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op72 (.out1(_69), .in1(ip_src_80_D), .in2(sbbit6_106_D));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op45 (.out1(_44), .in1(ip_dst_84_D), .in2(bsbit6_97_D));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op18 (.out1(_19), .in1(ip_dst_84_D), .in2(ssbit6_87_D));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op112 (.out1(R113), .clock(clock), .in1(_66));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op113 (.out1(R114), .clock(clock), .in1(_62));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op114 (.out1(R115), .clock(clock), .in1(_58));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op115 (.out1(R116), .clock(clock), .in1(_54));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op116 (.out1(R117), .clock(clock), .in1(_41));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op117 (.out1(R118), .clock(clock), .in1(_37));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op118 (.out1(R119), .clock(clock), .in1(_33));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op119 (.out1(R120), .clock(clock), .in1(_29));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op120 (.out1(R121), .clock(clock), .in1(_16));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op121 (.out1(R122), .clock(clock), .in1(_12));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op122 (.out1(R123), .clock(clock), .in1(_8));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op123 (.out1(R124), .clock(clock), .in1(_4));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op124 (.out1(R125), .clock(clock), .in1(_69));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op125 (.out1(R126), .clock(clock), .in1(_44));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op126 (.out1(R127), .clock(clock), .in1(_19));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(3), .BITSIZE_out1(32), .PRECISION(32)) op73 (.out1(_70), .in1(R125), .in2(3 'd 5));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(3), .BITSIZE_out1(32), .PRECISION(32)) op46 (.out1(_45), .in1(R126), .in2(3 'd 5));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(3), .BITSIZE_out1(32), .PRECISION(32)) op19 (.out1(_20), .in1(R127), .in2(3 'd 5));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op54 (.out1(_51), .in1(ip_src_80_D), .in2(sbbit1_101_D));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op27 (.out1(_26), .in1(ip_dst_84_D), .in2(bsbit1_92_D));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32), .PRECISION(32)) op0 (.out1(_1), .in1(ip_src_80_D), .in2(ssbit1_81_D));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(2), .BITSIZE_out1(32)) op58 (.out1(_55), .in1(R116), .in2(2 'd 2));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(1), .BITSIZE_out1(32)) op55 (.out1(_52), .in1(_51), .in2(1 'd 1));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(2), .BITSIZE_out1(32)) op31 (.out1(_30), .in1(R120), .in2(2 'd 2));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(1), .BITSIZE_out1(32)) op28 (.out1(_27), .in1(_26), .in2(1 'd 1));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(2), .BITSIZE_out1(32)) op4 (.out1(_5), .in1(R124), .in2(2 'd 2));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(1), .BITSIZE_out1(32)) op1 (.out1(_2), .in1(_1), .in2(1 'd 1));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(3), .BITSIZE_out1(32)) op62 (.out1(_59), .in1(R115), .in2(3 'd 4));
  bit_or #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op59 (.out1(_56), .in1(_52), .in2(_55));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(3), .BITSIZE_out1(32)) op35 (.out1(_34), .in1(R119), .in2(3 'd 4));
  bit_or #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op32 (.out1(_31), .in1(_27), .in2(_30));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(3), .BITSIZE_out1(32)) op8 (.out1(_9), .in1(R123), .in2(3 'd 4));
  bit_or #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op5 (.out1(_6), .in1(_2), .in2(_5));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(4), .BITSIZE_out1(32)) op66 (.out1(_63), .in1(R114), .in2(4 'd 8));
  bit_or #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op63 (.out1(_60), .in1(_56), .in2(_59));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(4), .BITSIZE_out1(32)) op39 (.out1(_38), .in1(R118), .in2(4 'd 8));
  bit_or #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op36 (.out1(_35), .in1(_31), .in2(_34));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(4), .BITSIZE_out1(32)) op12 (.out1(_13), .in1(R122), .in2(4 'd 8));
  bit_or #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op9 (.out1(_10), .in1(_6), .in2(_9));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(5), .BITSIZE_out1(32)) op70 (.out1(_67), .in1(R113), .in2(5 'd 16));
  bit_or #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op67 (.out1(_64), .in1(_60), .in2(_63));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(5), .BITSIZE_out1(32)) op43 (.out1(_42), .in1(R117), .in2(5 'd 16));
  bit_or #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op40 (.out1(_39), .in1(_35), .in2(_38));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(5), .BITSIZE_out1(32)) op16 (.out1(_17), .in1(R121), .in2(5 'd 16));
  bit_or #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op13 (.out1(_14), .in1(_10), .in2(_13));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op74 (.out1(_71), .in1(_70), .in2(6 'd 32));
  bit_or #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op71 (.out1(_68), .in1(_64), .in2(_67));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op47 (.out1(_46), .in1(_45), .in2(6 'd 32));
  bit_or #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op44 (.out1(_43), .in1(_39), .in2(_42));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op20 (.out1(_21), .in1(_20), .in2(6 'd 32));
  bit_or #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op17 (.out1(_18), .in1(_14), .in2(_17));
  bit_or #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op75 (.out1(_72), .in1(_68), .in2(_71));
  bit_or #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op48 (.out1(_47), .in1(_43), .in2(_46));
  bit_or #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op21 (.out1(_22), .in1(_18), .in2(_21));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op76 (.out1(sb_idx_107), .in1(_72));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op49 (.out1(bs_idx_98), .in1(_47));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op22 (.out1(ss_idx_88), .in1(_22));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op127 (.out1(R128), .clock(clock), .in1(sb_idx_107));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op128 (.out1(R129), .clock(clock), .in1(bs_idx_98));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op129 (.out1(R130), .clock(clock), .in1(ss_idx_88));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op77 (.out1(_73), .in1(R128));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op50 (.out1(_48), .in1(R129));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op23 (.out1(_23), .in1(R130));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op78 (.out1(_74), .in1(_73), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op51 (.out1(_49), .in1(_48), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op24 (.out1(_24), .in1(_23), .in2(2 'd 2));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op130 (.out1(R131), .clock(clock), .in1(_74));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op131 (.out1(R132), .clock(clock), .in1(_49));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op132 (.out1(R133), .clock(clock), .in1(_24));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op79 (.out1(_75), .in1(sb_subset_108_D), .in2(R131));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op52 (.out1(_50), .in1(bs_subset_99_D), .in2(R132));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op25 (.out1(_25), .in1(ss_subset_89_D), .in2(R133));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op133 (.out1(R134), .clock(clock), .in1(_75));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op134 (.out1(R135), .clock(clock), .in1(_50));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op135 (.out1(R136), .clock(clock), .in1(_25));
  SRAM op80 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(sb_leaf_109),.ADR(R134));
  SRAM op53 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(bs_leaf_100),.ADR(R135));
  SRAM op26 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(ss_leaf_91),.ADR(R136));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op136 (.out1(R137), .clock(clock), .in1(sb_leaf_109));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op137 (.out1(R138), .clock(clock), .in1(bs_leaf_100));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op138 (.out1(R139), .clock(clock), .in1(ss_leaf_91));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(5), .BITSIZE_out1(32), .PRECISION(32)) op88 (.out1(_78), .in1(R137), .in2(5 'd 16));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(5), .BITSIZE_out1(32), .PRECISION(32)) op85 (.out1(_77), .in1(R138), .in2(5 'd 16));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(5), .BITSIZE_out1(32), .PRECISION(32)) op82 (.out1(_76), .in1(R139), .in2(5 'd 16));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op84 (.out1(bs_priority_112), .in1(R138));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op81 (.out1(ss_priority_110), .in1(R139));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op87 (.out1(sb_priority_114), .in1(R137));
  GT_EXPR #(.BITSIZE_in1(16), .BITSIZE_in2(16),.BITSIZE_out1(1)) op90 (.out1(ifout90), .in1(ss_priority_110), .in2(bs_priority_112));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op89 (.out1(sb_matchid_115), .in1(_78));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op86 (.out1(bs_matchid_113), .in1(_77));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(16)) op83 (.out1(ss_matchid_111), .in1(_76));
  GT_EXPR #(.BITSIZE_in1(16), .BITSIZE_in2(16),.BITSIZE_out1(1)) op94 (.out1(ifout94), .in1(bs_priority_112), .in2(sb_priority_114));
  GT_EXPR #(.BITSIZE_in1(16), .BITSIZE_in2(16),.BITSIZE_out1(1)) op91 (.out1(ifout91), .in1(ss_priority_110), .in2(sb_priority_114));
  cast #(.BITSIZE_in1(16), .BITSIZE_out1(8)) op96 (.out1(_116), .in1(sb_matchid_115));
  cast #(.BITSIZE_in1(16), .BITSIZE_out1(8)) op95 (.out1(_117), .in1(bs_matchid_113));
  cast #(.BITSIZE_in1(16), .BITSIZE_out1(8)) op93 (.out1(_118), .in1(sb_matchid_115));
  cast #(.BITSIZE_in1(16), .BITSIZE_out1(8)) op92 (.out1(_119), .in1(ss_matchid_111));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op97 (.out1(mux0), .in1(_116), .in2(_117), .sel(ifout94));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op98 (.out1(mux1), .in1(_118), .in2(_119), .sel(ifout91));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op99 (.out1(mux2), .in1(mux0), .in2(mux1), .sel(ifout90));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op139 (.out1(R140), .clock(clock), .in1(mux2));
endmodule