`include "component_library.v"
`include "macros.v"

`timescale 1ns / 1ps
module top(clock, N16_233_D, N24_237_D, N32_241_D, N40_245_D, N48_249_D, N56_253_D, N64_257_D, N72_262_D, N80_266_D, N88_270_D, N96_274_D, N104_278_D, N112_282_D, N120_286_D, N128_289_D, C120_285_D, C112_281_D, C104_277_D, C96_273_D, C88_269_D, C80_265_D, C72_261_D, ip2_259_D, C64_256_D, C56_252_D, C48_248_D, C40_244_D, C32_240_D, C24_236_D, C16_231_D, ip1_229_D, R2336);
  //IN
  input clock;
  input [63:0] N16_233_D;
  input [63:0] N24_237_D;
  input [63:0] N32_241_D;
  input [63:0] N40_245_D;
  input [63:0] N48_249_D;
  input [63:0] N56_253_D;
  input [63:0] N64_257_D;
  input [63:0] N72_262_D;
  input [63:0] N80_266_D;
  input [63:0] N88_270_D;
  input [63:0] N96_274_D;
  input [63:0] N104_278_D;
  input [63:0] N112_282_D;
  input [63:0] N120_286_D;
  input [63:0] N128_289_D;
  input [63:0] C120_285_D;
  input [63:0] C112_281_D;
  input [63:0] C104_277_D;
  input [63:0] C96_273_D;
  input [63:0] C88_269_D;
  input [63:0] C80_265_D;
  input [63:0] C72_261_D;
  input [63:0] ip2_259_D;
  input [63:0] C64_256_D;
  input [63:0] C56_252_D;
  input [63:0] C48_248_D;
  input [63:0] C40_244_D;
  input [63:0] C32_240_D;
  input [63:0] C24_236_D;
  input [63:0] C16_231_D;
  input [63:0] ip1_229_D;
  //OUT
  output [7:0] R2336;
  //WIRES
  wire [7:0] R2336;
  wire [7:0] R2335;
  wire [7:0] R2334;
  wire [7:0] R2333;
  wire [7:0] R2332;
  wire [7:0] R2331;
  wire [7:0] R2330;
  wire [7:0] R2329;
  wire [7:0] R2328;
  wire [7:0] R2327;
  wire [63:0] R2326;
  wire [63:0] R2325;
  wire [63:0] R2324;
  wire [63:0] R2323;
  wire [63:0] R2322;
  wire [63:0] R2321;
  wire [7:0] R2320;
  wire [7:0] R2319;
  wire [7:0] R2318;
  wire [7:0] R2317;
  wire [7:0] R2316;
  wire [7:0] R2315;
  wire [7:0] R2314;
  wire [7:0] R2313;
  wire [7:0] R2312;
  wire [63:0] R2311;
  wire [63:0] R2310;
  wire [63:0] R2309;
  wire [63:0] R2308;
  wire [63:0] R2307;
  wire [63:0] R2306;
  wire [63:0] R2305;
  wire [63:0] R2304;
  wire [63:0] R2303;
  wire [31:0] R2302;
  wire [31:0] R2301;
  wire [31:0] R2300;
  wire [31:0] R2299;
  wire [63:0] R2298;
  wire [63:0] R2297;
  wire [0:0] R2296;
  wire [0:0] R2295;
  wire [0:0] R2294;
  wire [0:0] R2293;
  wire [0:0] R2292;
  wire [0:0] R2291;
  wire [0:0] R2290;
  wire [0:0] R2289;
  wire [31:0] R2288;
  wire [63:0] R2287;
  wire [63:0] R2286;
  wire [31:0] R2285;
  wire [31:0] R2284;
  wire [31:0] R2283;
  wire [31:0] R2282;
  wire [31:0] R2281;
  wire [31:0] R2280;
  wire [31:0] R2279;
  wire [31:0] R2278;
  wire [31:0] R2277;
  wire [31:0] R2276;
  wire [31:0] R2275;
  wire [31:0] R2274;
  wire [31:0] R2273;
  wire [63:0] R2272;
  wire [63:0] R2271;
  wire [0:0] R2270;
  wire [0:0] R2269;
  wire [0:0] R2268;
  wire [0:0] R2267;
  wire [0:0] R2266;
  wire [0:0] R2265;
  wire [0:0] R2264;
  wire [0:0] R2263;
  wire [0:0] R2262;
  wire [0:0] R2261;
  wire [0:0] R2260;
  wire [0:0] R2259;
  wire [0:0] R2258;
  wire [0:0] R2257;
  wire [0:0] R2256;
  wire [0:0] R2255;
  wire [0:0] R2254;
  wire [31:0] R2253;
  wire [63:0] R2252;
  wire [63:0] R2251;
  wire [31:0] R2250;
  wire [31:0] R2249;
  wire [31:0] R2248;
  wire [31:0] R2247;
  wire [31:0] R2246;
  wire [31:0] R2245;
  wire [31:0] R2244;
  wire [31:0] R2243;
  wire [31:0] R2242;
  wire [31:0] R2241;
  wire [31:0] R2240;
  wire [31:0] R2239;
  wire [31:0] R2238;
  wire [31:0] R2237;
  wire [31:0] R2236;
  wire [31:0] R2235;
  wire [31:0] R2234;
  wire [31:0] R2233;
  wire [31:0] R2232;
  wire [31:0] R2231;
  wire [31:0] R2230;
  wire [31:0] R2229;
  wire [63:0] R2228;
  wire [63:0] R2227;
  wire [0:0] R2226;
  wire [0:0] R2225;
  wire [0:0] R2224;
  wire [0:0] R2223;
  wire [0:0] R2222;
  wire [0:0] R2221;
  wire [0:0] R2220;
  wire [0:0] R2219;
  wire [0:0] R2218;
  wire [0:0] R2217;
  wire [0:0] R2216;
  wire [0:0] R2215;
  wire [0:0] R2214;
  wire [0:0] R2213;
  wire [0:0] R2212;
  wire [0:0] R2211;
  wire [0:0] R2210;
  wire [0:0] R2209;
  wire [0:0] R2208;
  wire [0:0] R2207;
  wire [0:0] R2206;
  wire [0:0] R2205;
  wire [0:0] R2204;
  wire [0:0] R2203;
  wire [0:0] R2202;
  wire [0:0] R2201;
  wire [31:0] R2200;
  wire [63:0] R2199;
  wire [63:0] R2198;
  wire [31:0] R2197;
  wire [31:0] R2196;
  wire [31:0] R2195;
  wire [31:0] R2194;
  wire [31:0] R2193;
  wire [31:0] R2192;
  wire [31:0] R2191;
  wire [31:0] R2190;
  wire [31:0] R2189;
  wire [31:0] R2188;
  wire [31:0] R2187;
  wire [31:0] R2186;
  wire [31:0] R2185;
  wire [31:0] R2184;
  wire [31:0] R2183;
  wire [31:0] R2182;
  wire [31:0] R2181;
  wire [31:0] R2180;
  wire [31:0] R2179;
  wire [31:0] R2178;
  wire [31:0] R2177;
  wire [31:0] R2176;
  wire [31:0] R2175;
  wire [31:0] R2174;
  wire [31:0] R2173;
  wire [31:0] R2172;
  wire [31:0] R2171;
  wire [31:0] R2170;
  wire [31:0] R2169;
  wire [31:0] R2168;
  wire [31:0] R2167;
  wire [63:0] R2166;
  wire [63:0] R2165;
  wire [0:0] R2164;
  wire [0:0] R2163;
  wire [0:0] R2162;
  wire [0:0] R2161;
  wire [0:0] R2160;
  wire [0:0] R2159;
  wire [0:0] R2158;
  wire [0:0] R2157;
  wire [0:0] R2156;
  wire [0:0] R2155;
  wire [0:0] R2154;
  wire [0:0] R2153;
  wire [0:0] R2152;
  wire [0:0] R2151;
  wire [0:0] R2150;
  wire [0:0] R2149;
  wire [0:0] R2148;
  wire [0:0] R2147;
  wire [0:0] R2146;
  wire [0:0] R2145;
  wire [0:0] R2144;
  wire [0:0] R2143;
  wire [0:0] R2142;
  wire [0:0] R2141;
  wire [0:0] R2140;
  wire [0:0] R2139;
  wire [0:0] R2138;
  wire [0:0] R2137;
  wire [0:0] R2136;
  wire [0:0] R2135;
  wire [0:0] R2134;
  wire [0:0] R2133;
  wire [0:0] R2132;
  wire [0:0] R2131;
  wire [0:0] R2130;
  wire [31:0] R2129;
  wire [63:0] R2128;
  wire [63:0] R2127;
  wire [31:0] R2126;
  wire [31:0] R2125;
  wire [31:0] R2124;
  wire [31:0] R2123;
  wire [31:0] R2122;
  wire [31:0] R2121;
  wire [31:0] R2120;
  wire [31:0] R2119;
  wire [31:0] R2118;
  wire [31:0] R2117;
  wire [31:0] R2116;
  wire [31:0] R2115;
  wire [31:0] R2114;
  wire [31:0] R2113;
  wire [31:0] R2112;
  wire [31:0] R2111;
  wire [31:0] R2110;
  wire [31:0] R2109;
  wire [31:0] R2108;
  wire [31:0] R2107;
  wire [31:0] R2106;
  wire [31:0] R2105;
  wire [31:0] R2104;
  wire [31:0] R2103;
  wire [31:0] R2102;
  wire [31:0] R2101;
  wire [31:0] R2100;
  wire [31:0] R2099;
  wire [31:0] R2098;
  wire [31:0] R2097;
  wire [31:0] R2096;
  wire [31:0] R2095;
  wire [31:0] R2094;
  wire [31:0] R2093;
  wire [31:0] R2092;
  wire [31:0] R2091;
  wire [31:0] R2090;
  wire [31:0] R2089;
  wire [31:0] R2088;
  wire [31:0] R2087;
  wire [63:0] R2086;
  wire [63:0] R2085;
  wire [0:0] R2084;
  wire [0:0] R2083;
  wire [0:0] R2082;
  wire [0:0] R2081;
  wire [0:0] R2080;
  wire [0:0] R2079;
  wire [0:0] R2078;
  wire [0:0] R2077;
  wire [0:0] R2076;
  wire [0:0] R2075;
  wire [0:0] R2074;
  wire [0:0] R2073;
  wire [0:0] R2072;
  wire [0:0] R2071;
  wire [0:0] R2070;
  wire [0:0] R2069;
  wire [0:0] R2068;
  wire [0:0] R2067;
  wire [0:0] R2066;
  wire [0:0] R2065;
  wire [0:0] R2064;
  wire [0:0] R2063;
  wire [0:0] R2062;
  wire [0:0] R2061;
  wire [0:0] R2060;
  wire [0:0] R2059;
  wire [0:0] R2058;
  wire [0:0] R2057;
  wire [0:0] R2056;
  wire [0:0] R2055;
  wire [0:0] R2054;
  wire [0:0] R2053;
  wire [0:0] R2052;
  wire [0:0] R2051;
  wire [0:0] R2050;
  wire [0:0] R2049;
  wire [0:0] R2048;
  wire [0:0] R2047;
  wire [0:0] R2046;
  wire [0:0] R2045;
  wire [0:0] R2044;
  wire [0:0] R2043;
  wire [0:0] R2042;
  wire [0:0] R2041;
  wire [31:0] R2040;
  wire [63:0] R2039;
  wire [63:0] R2038;
  wire [31:0] R2037;
  wire [31:0] R2036;
  wire [31:0] R2035;
  wire [31:0] R2034;
  wire [31:0] R2033;
  wire [31:0] R2032;
  wire [31:0] R2031;
  wire [31:0] R2030;
  wire [31:0] R2029;
  wire [31:0] R2028;
  wire [31:0] R2027;
  wire [31:0] R2026;
  wire [31:0] R2025;
  wire [31:0] R2024;
  wire [31:0] R2023;
  wire [31:0] R2022;
  wire [31:0] R2021;
  wire [31:0] R2020;
  wire [31:0] R2019;
  wire [31:0] R2018;
  wire [31:0] R2017;
  wire [31:0] R2016;
  wire [31:0] R2015;
  wire [31:0] R2014;
  wire [31:0] R2013;
  wire [31:0] R2012;
  wire [31:0] R2011;
  wire [31:0] R2010;
  wire [31:0] R2009;
  wire [31:0] R2008;
  wire [31:0] R2007;
  wire [31:0] R2006;
  wire [31:0] R2005;
  wire [31:0] R2004;
  wire [31:0] R2003;
  wire [31:0] R2002;
  wire [31:0] R2001;
  wire [31:0] R2000;
  wire [31:0] R1999;
  wire [31:0] R1998;
  wire [31:0] R1997;
  wire [31:0] R1996;
  wire [31:0] R1995;
  wire [31:0] R1994;
  wire [31:0] R1993;
  wire [31:0] R1992;
  wire [31:0] R1991;
  wire [31:0] R1990;
  wire [31:0] R1989;
  wire [63:0] R1988;
  wire [63:0] R1987;
  wire [0:0] R1986;
  wire [0:0] R1985;
  wire [0:0] R1984;
  wire [0:0] R1983;
  wire [0:0] R1982;
  wire [0:0] R1981;
  wire [0:0] R1980;
  wire [0:0] R1979;
  wire [0:0] R1978;
  wire [0:0] R1977;
  wire [0:0] R1976;
  wire [0:0] R1975;
  wire [0:0] R1974;
  wire [0:0] R1973;
  wire [0:0] R1972;
  wire [0:0] R1971;
  wire [0:0] R1970;
  wire [0:0] R1969;
  wire [0:0] R1968;
  wire [0:0] R1967;
  wire [0:0] R1966;
  wire [0:0] R1965;
  wire [0:0] R1964;
  wire [0:0] R1963;
  wire [0:0] R1962;
  wire [0:0] R1961;
  wire [0:0] R1960;
  wire [0:0] R1959;
  wire [0:0] R1958;
  wire [0:0] R1957;
  wire [0:0] R1956;
  wire [0:0] R1955;
  wire [0:0] R1954;
  wire [0:0] R1953;
  wire [0:0] R1952;
  wire [0:0] R1951;
  wire [0:0] R1950;
  wire [0:0] R1949;
  wire [0:0] R1948;
  wire [0:0] R1947;
  wire [0:0] R1946;
  wire [0:0] R1945;
  wire [0:0] R1944;
  wire [0:0] R1943;
  wire [0:0] R1942;
  wire [0:0] R1941;
  wire [0:0] R1940;
  wire [0:0] R1939;
  wire [0:0] R1938;
  wire [0:0] R1937;
  wire [0:0] R1936;
  wire [0:0] R1935;
  wire [0:0] R1934;
  wire [31:0] R1933;
  wire [63:0] R1932;
  wire [63:0] R1931;
  wire [31:0] R1930;
  wire [31:0] R1929;
  wire [31:0] R1928;
  wire [31:0] R1927;
  wire [31:0] R1926;
  wire [31:0] R1925;
  wire [31:0] R1924;
  wire [31:0] R1923;
  wire [31:0] R1922;
  wire [31:0] R1921;
  wire [31:0] R1920;
  wire [31:0] R1919;
  wire [31:0] R1918;
  wire [31:0] R1917;
  wire [31:0] R1916;
  wire [31:0] R1915;
  wire [31:0] R1914;
  wire [31:0] R1913;
  wire [31:0] R1912;
  wire [31:0] R1911;
  wire [31:0] R1910;
  wire [31:0] R1909;
  wire [31:0] R1908;
  wire [31:0] R1907;
  wire [31:0] R1906;
  wire [31:0] R1905;
  wire [31:0] R1904;
  wire [31:0] R1903;
  wire [31:0] R1902;
  wire [31:0] R1901;
  wire [31:0] R1900;
  wire [31:0] R1899;
  wire [31:0] R1898;
  wire [31:0] R1897;
  wire [31:0] R1896;
  wire [31:0] R1895;
  wire [31:0] R1894;
  wire [31:0] R1893;
  wire [31:0] R1892;
  wire [31:0] R1891;
  wire [31:0] R1890;
  wire [31:0] R1889;
  wire [31:0] R1888;
  wire [31:0] R1887;
  wire [31:0] R1886;
  wire [31:0] R1885;
  wire [31:0] R1884;
  wire [31:0] R1883;
  wire [31:0] R1882;
  wire [31:0] R1881;
  wire [31:0] R1880;
  wire [31:0] R1879;
  wire [31:0] R1878;
  wire [31:0] R1877;
  wire [31:0] R1876;
  wire [31:0] R1875;
  wire [31:0] R1874;
  wire [31:0] R1873;
  wire [63:0] R1872;
  wire [63:0] R1871;
  wire [0:0] R1870;
  wire [0:0] R1869;
  wire [0:0] R1868;
  wire [0:0] R1867;
  wire [0:0] R1866;
  wire [0:0] R1865;
  wire [0:0] R1864;
  wire [0:0] R1863;
  wire [0:0] R1862;
  wire [0:0] R1861;
  wire [0:0] R1860;
  wire [0:0] R1859;
  wire [0:0] R1858;
  wire [0:0] R1857;
  wire [0:0] R1856;
  wire [0:0] R1855;
  wire [0:0] R1854;
  wire [0:0] R1853;
  wire [0:0] R1852;
  wire [0:0] R1851;
  wire [0:0] R1850;
  wire [0:0] R1849;
  wire [0:0] R1848;
  wire [0:0] R1847;
  wire [0:0] R1846;
  wire [0:0] R1845;
  wire [0:0] R1844;
  wire [0:0] R1843;
  wire [0:0] R1842;
  wire [0:0] R1841;
  wire [0:0] R1840;
  wire [0:0] R1839;
  wire [0:0] R1838;
  wire [0:0] R1837;
  wire [0:0] R1836;
  wire [0:0] R1835;
  wire [0:0] R1834;
  wire [0:0] R1833;
  wire [0:0] R1832;
  wire [0:0] R1831;
  wire [0:0] R1830;
  wire [0:0] R1829;
  wire [0:0] R1828;
  wire [0:0] R1827;
  wire [0:0] R1826;
  wire [0:0] R1825;
  wire [0:0] R1824;
  wire [0:0] R1823;
  wire [0:0] R1822;
  wire [0:0] R1821;
  wire [0:0] R1820;
  wire [0:0] R1819;
  wire [0:0] R1818;
  wire [0:0] R1817;
  wire [0:0] R1816;
  wire [0:0] R1815;
  wire [0:0] R1814;
  wire [0:0] R1813;
  wire [0:0] R1812;
  wire [0:0] R1811;
  wire [0:0] R1810;
  wire [0:0] R1809;
  wire [0:0] R1808;
  wire [31:0] R1807;
  wire [63:0] R1806;
  wire [63:0] R1805;
  wire [31:0] R1804;
  wire [31:0] R1803;
  wire [31:0] R1802;
  wire [31:0] R1801;
  wire [31:0] R1800;
  wire [31:0] R1799;
  wire [31:0] R1798;
  wire [31:0] R1797;
  wire [31:0] R1796;
  wire [31:0] R1795;
  wire [31:0] R1794;
  wire [31:0] R1793;
  wire [31:0] R1792;
  wire [31:0] R1791;
  wire [31:0] R1790;
  wire [31:0] R1789;
  wire [31:0] R1788;
  wire [31:0] R1787;
  wire [31:0] R1786;
  wire [31:0] R1785;
  wire [31:0] R1784;
  wire [31:0] R1783;
  wire [31:0] R1782;
  wire [31:0] R1781;
  wire [31:0] R1780;
  wire [31:0] R1779;
  wire [31:0] R1778;
  wire [31:0] R1777;
  wire [31:0] R1776;
  wire [31:0] R1775;
  wire [31:0] R1774;
  wire [31:0] R1773;
  wire [31:0] R1772;
  wire [31:0] R1771;
  wire [31:0] R1770;
  wire [31:0] R1769;
  wire [31:0] R1768;
  wire [31:0] R1767;
  wire [31:0] R1766;
  wire [31:0] R1765;
  wire [31:0] R1764;
  wire [31:0] R1763;
  wire [31:0] R1762;
  wire [31:0] R1761;
  wire [31:0] R1760;
  wire [31:0] R1759;
  wire [31:0] R1758;
  wire [31:0] R1757;
  wire [31:0] R1756;
  wire [31:0] R1755;
  wire [31:0] R1754;
  wire [31:0] R1753;
  wire [31:0] R1752;
  wire [31:0] R1751;
  wire [31:0] R1750;
  wire [31:0] R1749;
  wire [31:0] R1748;
  wire [31:0] R1747;
  wire [31:0] R1746;
  wire [31:0] R1745;
  wire [31:0] R1744;
  wire [31:0] R1743;
  wire [31:0] R1742;
  wire [31:0] R1741;
  wire [31:0] R1740;
  wire [31:0] R1739;
  wire [31:0] R1738;
  wire [63:0] R1737;
  wire [63:0] R1736;
  wire [0:0] R1735;
  wire [0:0] R1734;
  wire [0:0] R1733;
  wire [0:0] R1732;
  wire [0:0] R1731;
  wire [0:0] R1730;
  wire [0:0] R1729;
  wire [0:0] R1728;
  wire [0:0] R1727;
  wire [0:0] R1726;
  wire [0:0] R1725;
  wire [0:0] R1724;
  wire [0:0] R1723;
  wire [0:0] R1722;
  wire [0:0] R1721;
  wire [0:0] R1720;
  wire [0:0] R1719;
  wire [0:0] R1718;
  wire [0:0] R1717;
  wire [0:0] R1716;
  wire [0:0] R1715;
  wire [0:0] R1714;
  wire [0:0] R1713;
  wire [0:0] R1712;
  wire [0:0] R1711;
  wire [0:0] R1710;
  wire [0:0] R1709;
  wire [0:0] R1708;
  wire [0:0] R1707;
  wire [0:0] R1706;
  wire [0:0] R1705;
  wire [0:0] R1704;
  wire [0:0] R1703;
  wire [0:0] R1702;
  wire [0:0] R1701;
  wire [0:0] R1700;
  wire [0:0] R1699;
  wire [0:0] R1698;
  wire [0:0] R1697;
  wire [0:0] R1696;
  wire [0:0] R1695;
  wire [0:0] R1694;
  wire [0:0] R1693;
  wire [0:0] R1692;
  wire [0:0] R1691;
  wire [0:0] R1690;
  wire [0:0] R1689;
  wire [0:0] R1688;
  wire [0:0] R1687;
  wire [0:0] R1686;
  wire [0:0] R1685;
  wire [0:0] R1684;
  wire [0:0] R1683;
  wire [0:0] R1682;
  wire [0:0] R1681;
  wire [0:0] R1680;
  wire [0:0] R1679;
  wire [0:0] R1678;
  wire [0:0] R1677;
  wire [0:0] R1676;
  wire [0:0] R1675;
  wire [0:0] R1674;
  wire [0:0] R1673;
  wire [0:0] R1672;
  wire [0:0] R1671;
  wire [0:0] R1670;
  wire [0:0] R1669;
  wire [0:0] R1668;
  wire [0:0] R1667;
  wire [0:0] R1666;
  wire [0:0] R1665;
  wire [0:0] R1664;
  wire [31:0] R1663;
  wire [63:0] R1662;
  wire [63:0] R1661;
  wire [31:0] R1660;
  wire [31:0] R1659;
  wire [31:0] R1658;
  wire [31:0] R1657;
  wire [31:0] R1656;
  wire [31:0] R1655;
  wire [31:0] R1654;
  wire [31:0] R1653;
  wire [31:0] R1652;
  wire [31:0] R1651;
  wire [31:0] R1650;
  wire [31:0] R1649;
  wire [31:0] R1648;
  wire [31:0] R1647;
  wire [31:0] R1646;
  wire [31:0] R1645;
  wire [31:0] R1644;
  wire [31:0] R1643;
  wire [31:0] R1642;
  wire [31:0] R1641;
  wire [31:0] R1640;
  wire [31:0] R1639;
  wire [31:0] R1638;
  wire [31:0] R1637;
  wire [31:0] R1636;
  wire [31:0] R1635;
  wire [31:0] R1634;
  wire [31:0] R1633;
  wire [31:0] R1632;
  wire [31:0] R1631;
  wire [31:0] R1630;
  wire [31:0] R1629;
  wire [31:0] R1628;
  wire [31:0] R1627;
  wire [31:0] R1626;
  wire [31:0] R1625;
  wire [31:0] R1624;
  wire [31:0] R1623;
  wire [31:0] R1622;
  wire [31:0] R1621;
  wire [31:0] R1620;
  wire [31:0] R1619;
  wire [31:0] R1618;
  wire [31:0] R1617;
  wire [31:0] R1616;
  wire [31:0] R1615;
  wire [31:0] R1614;
  wire [31:0] R1613;
  wire [31:0] R1612;
  wire [31:0] R1611;
  wire [31:0] R1610;
  wire [31:0] R1609;
  wire [31:0] R1608;
  wire [31:0] R1607;
  wire [31:0] R1606;
  wire [31:0] R1605;
  wire [31:0] R1604;
  wire [31:0] R1603;
  wire [31:0] R1602;
  wire [31:0] R1601;
  wire [31:0] R1600;
  wire [31:0] R1599;
  wire [31:0] R1598;
  wire [31:0] R1597;
  wire [31:0] R1596;
  wire [31:0] R1595;
  wire [31:0] R1594;
  wire [31:0] R1593;
  wire [31:0] R1592;
  wire [31:0] R1591;
  wire [31:0] R1590;
  wire [31:0] R1589;
  wire [31:0] R1588;
  wire [31:0] R1587;
  wire [31:0] R1586;
  wire [31:0] R1585;
  wire [63:0] R1584;
  wire [63:0] R1583;
  wire [0:0] R1582;
  wire [0:0] R1581;
  wire [0:0] R1580;
  wire [0:0] R1579;
  wire [0:0] R1578;
  wire [0:0] R1577;
  wire [0:0] R1576;
  wire [0:0] R1575;
  wire [0:0] R1574;
  wire [0:0] R1573;
  wire [0:0] R1572;
  wire [0:0] R1571;
  wire [0:0] R1570;
  wire [0:0] R1569;
  wire [0:0] R1568;
  wire [0:0] R1567;
  wire [0:0] R1566;
  wire [0:0] R1565;
  wire [0:0] R1564;
  wire [0:0] R1563;
  wire [0:0] R1562;
  wire [0:0] R1561;
  wire [0:0] R1560;
  wire [0:0] R1559;
  wire [0:0] R1558;
  wire [0:0] R1557;
  wire [0:0] R1556;
  wire [0:0] R1555;
  wire [0:0] R1554;
  wire [0:0] R1553;
  wire [0:0] R1552;
  wire [0:0] R1551;
  wire [0:0] R1550;
  wire [0:0] R1549;
  wire [0:0] R1548;
  wire [0:0] R1547;
  wire [0:0] R1546;
  wire [0:0] R1545;
  wire [0:0] R1544;
  wire [0:0] R1543;
  wire [0:0] R1542;
  wire [0:0] R1541;
  wire [0:0] R1540;
  wire [0:0] R1539;
  wire [0:0] R1538;
  wire [0:0] R1537;
  wire [0:0] R1536;
  wire [0:0] R1535;
  wire [0:0] R1534;
  wire [0:0] R1533;
  wire [0:0] R1532;
  wire [0:0] R1531;
  wire [0:0] R1530;
  wire [0:0] R1529;
  wire [0:0] R1528;
  wire [0:0] R1527;
  wire [0:0] R1526;
  wire [0:0] R1525;
  wire [0:0] R1524;
  wire [0:0] R1523;
  wire [0:0] R1522;
  wire [0:0] R1521;
  wire [0:0] R1520;
  wire [0:0] R1519;
  wire [0:0] R1518;
  wire [0:0] R1517;
  wire [0:0] R1516;
  wire [0:0] R1515;
  wire [0:0] R1514;
  wire [0:0] R1513;
  wire [0:0] R1512;
  wire [0:0] R1511;
  wire [0:0] R1510;
  wire [0:0] R1509;
  wire [0:0] R1508;
  wire [0:0] R1507;
  wire [0:0] R1506;
  wire [0:0] R1505;
  wire [0:0] R1504;
  wire [0:0] R1503;
  wire [0:0] R1502;
  wire [31:0] R1501;
  wire [63:0] R1500;
  wire [63:0] R1499;
  wire [31:0] R1498;
  wire [31:0] R1497;
  wire [31:0] R1496;
  wire [31:0] R1495;
  wire [31:0] R1494;
  wire [31:0] R1493;
  wire [31:0] R1492;
  wire [31:0] R1491;
  wire [31:0] R1490;
  wire [31:0] R1489;
  wire [31:0] R1488;
  wire [31:0] R1487;
  wire [31:0] R1486;
  wire [31:0] R1485;
  wire [31:0] R1484;
  wire [31:0] R1483;
  wire [31:0] R1482;
  wire [31:0] R1481;
  wire [31:0] R1480;
  wire [31:0] R1479;
  wire [31:0] R1478;
  wire [31:0] R1477;
  wire [31:0] R1476;
  wire [31:0] R1475;
  wire [31:0] R1474;
  wire [31:0] R1473;
  wire [31:0] R1472;
  wire [31:0] R1471;
  wire [31:0] R1470;
  wire [31:0] R1469;
  wire [31:0] R1468;
  wire [31:0] R1467;
  wire [31:0] R1466;
  wire [31:0] R1465;
  wire [31:0] R1464;
  wire [31:0] R1463;
  wire [31:0] R1462;
  wire [31:0] R1461;
  wire [31:0] R1460;
  wire [31:0] R1459;
  wire [31:0] R1458;
  wire [31:0] R1457;
  wire [31:0] R1456;
  wire [31:0] R1455;
  wire [31:0] R1454;
  wire [31:0] R1453;
  wire [31:0] R1452;
  wire [31:0] R1451;
  wire [31:0] R1450;
  wire [31:0] R1449;
  wire [31:0] R1448;
  wire [31:0] R1447;
  wire [31:0] R1446;
  wire [31:0] R1445;
  wire [31:0] R1444;
  wire [31:0] R1443;
  wire [31:0] R1442;
  wire [31:0] R1441;
  wire [31:0] R1440;
  wire [31:0] R1439;
  wire [31:0] R1438;
  wire [31:0] R1437;
  wire [31:0] R1436;
  wire [31:0] R1435;
  wire [31:0] R1434;
  wire [31:0] R1433;
  wire [31:0] R1432;
  wire [31:0] R1431;
  wire [31:0] R1430;
  wire [31:0] R1429;
  wire [31:0] R1428;
  wire [31:0] R1427;
  wire [31:0] R1426;
  wire [31:0] R1425;
  wire [31:0] R1424;
  wire [31:0] R1423;
  wire [31:0] R1422;
  wire [31:0] R1421;
  wire [31:0] R1420;
  wire [31:0] R1419;
  wire [31:0] R1418;
  wire [31:0] R1417;
  wire [31:0] R1416;
  wire [31:0] R1415;
  wire [31:0] R1414;
  wire [31:0] R1413;
  wire [63:0] R1412;
  wire [63:0] R1411;
  wire [0:0] R1410;
  wire [0:0] R1409;
  wire [0:0] R1408;
  wire [0:0] R1407;
  wire [0:0] R1406;
  wire [0:0] R1405;
  wire [0:0] R1404;
  wire [0:0] R1403;
  wire [0:0] R1402;
  wire [0:0] R1401;
  wire [0:0] R1400;
  wire [0:0] R1399;
  wire [0:0] R1398;
  wire [0:0] R1397;
  wire [0:0] R1396;
  wire [0:0] R1395;
  wire [0:0] R1394;
  wire [0:0] R1393;
  wire [0:0] R1392;
  wire [0:0] R1391;
  wire [0:0] R1390;
  wire [0:0] R1389;
  wire [0:0] R1388;
  wire [0:0] R1387;
  wire [0:0] R1386;
  wire [0:0] R1385;
  wire [0:0] R1384;
  wire [0:0] R1383;
  wire [0:0] R1382;
  wire [0:0] R1381;
  wire [0:0] R1380;
  wire [0:0] R1379;
  wire [0:0] R1378;
  wire [0:0] R1377;
  wire [0:0] R1376;
  wire [0:0] R1375;
  wire [0:0] R1374;
  wire [0:0] R1373;
  wire [0:0] R1372;
  wire [0:0] R1371;
  wire [0:0] R1370;
  wire [0:0] R1369;
  wire [0:0] R1368;
  wire [0:0] R1367;
  wire [0:0] R1366;
  wire [0:0] R1365;
  wire [0:0] R1364;
  wire [0:0] R1363;
  wire [0:0] R1362;
  wire [0:0] R1361;
  wire [0:0] R1360;
  wire [0:0] R1359;
  wire [0:0] R1358;
  wire [0:0] R1357;
  wire [0:0] R1356;
  wire [0:0] R1355;
  wire [0:0] R1354;
  wire [0:0] R1353;
  wire [0:0] R1352;
  wire [0:0] R1351;
  wire [0:0] R1350;
  wire [0:0] R1349;
  wire [0:0] R1348;
  wire [0:0] R1347;
  wire [0:0] R1346;
  wire [0:0] R1345;
  wire [0:0] R1344;
  wire [0:0] R1343;
  wire [0:0] R1342;
  wire [0:0] R1341;
  wire [0:0] R1340;
  wire [0:0] R1339;
  wire [0:0] R1338;
  wire [0:0] R1337;
  wire [0:0] R1336;
  wire [0:0] R1335;
  wire [0:0] R1334;
  wire [0:0] R1333;
  wire [0:0] R1332;
  wire [0:0] R1331;
  wire [0:0] R1330;
  wire [0:0] R1329;
  wire [0:0] R1328;
  wire [0:0] R1327;
  wire [0:0] R1326;
  wire [0:0] R1325;
  wire [0:0] R1324;
  wire [0:0] R1323;
  wire [0:0] R1322;
  wire [0:0] R1321;
  wire [31:0] R1320;
  wire [63:0] R1319;
  wire [63:0] R1318;
  wire [31:0] R1317;
  wire [31:0] R1316;
  wire [31:0] R1315;
  wire [31:0] R1314;
  wire [31:0] R1313;
  wire [31:0] R1312;
  wire [31:0] R1311;
  wire [31:0] R1310;
  wire [31:0] R1309;
  wire [31:0] R1308;
  wire [31:0] R1307;
  wire [31:0] R1306;
  wire [31:0] R1305;
  wire [31:0] R1304;
  wire [31:0] R1303;
  wire [31:0] R1302;
  wire [31:0] R1301;
  wire [31:0] R1300;
  wire [31:0] R1299;
  wire [31:0] R1298;
  wire [31:0] R1297;
  wire [31:0] R1296;
  wire [31:0] R1295;
  wire [31:0] R1294;
  wire [31:0] R1293;
  wire [31:0] R1292;
  wire [31:0] R1291;
  wire [31:0] R1290;
  wire [31:0] R1289;
  wire [31:0] R1288;
  wire [31:0] R1287;
  wire [31:0] R1286;
  wire [31:0] R1285;
  wire [31:0] R1284;
  wire [31:0] R1283;
  wire [31:0] R1282;
  wire [31:0] R1281;
  wire [31:0] R1280;
  wire [31:0] R1279;
  wire [31:0] R1278;
  wire [31:0] R1277;
  wire [31:0] R1276;
  wire [31:0] R1275;
  wire [31:0] R1274;
  wire [31:0] R1273;
  wire [31:0] R1272;
  wire [31:0] R1271;
  wire [31:0] R1270;
  wire [31:0] R1269;
  wire [31:0] R1268;
  wire [31:0] R1267;
  wire [31:0] R1266;
  wire [31:0] R1265;
  wire [31:0] R1264;
  wire [31:0] R1263;
  wire [31:0] R1262;
  wire [31:0] R1261;
  wire [31:0] R1260;
  wire [31:0] R1259;
  wire [31:0] R1258;
  wire [31:0] R1257;
  wire [31:0] R1256;
  wire [31:0] R1255;
  wire [31:0] R1254;
  wire [31:0] R1253;
  wire [31:0] R1252;
  wire [31:0] R1251;
  wire [31:0] R1250;
  wire [31:0] R1249;
  wire [31:0] R1248;
  wire [31:0] R1247;
  wire [31:0] R1246;
  wire [31:0] R1245;
  wire [31:0] R1244;
  wire [31:0] R1243;
  wire [31:0] R1242;
  wire [31:0] R1241;
  wire [31:0] R1240;
  wire [31:0] R1239;
  wire [31:0] R1238;
  wire [31:0] R1237;
  wire [31:0] R1236;
  wire [31:0] R1235;
  wire [31:0] R1234;
  wire [31:0] R1233;
  wire [31:0] R1232;
  wire [31:0] R1231;
  wire [31:0] R1230;
  wire [31:0] R1229;
  wire [31:0] R1228;
  wire [31:0] R1227;
  wire [31:0] R1226;
  wire [31:0] R1225;
  wire [31:0] R1224;
  wire [31:0] R1223;
  wire [63:0] R1222;
  wire [63:0] R1221;
  wire [0:0] R1220;
  wire [0:0] R1219;
  wire [0:0] R1218;
  wire [0:0] R1217;
  wire [0:0] R1216;
  wire [0:0] R1215;
  wire [0:0] R1214;
  wire [0:0] R1213;
  wire [0:0] R1212;
  wire [0:0] R1211;
  wire [0:0] R1210;
  wire [0:0] R1209;
  wire [0:0] R1208;
  wire [0:0] R1207;
  wire [0:0] R1206;
  wire [0:0] R1205;
  wire [0:0] R1204;
  wire [0:0] R1203;
  wire [0:0] R1202;
  wire [0:0] R1201;
  wire [0:0] R1200;
  wire [0:0] R1199;
  wire [0:0] R1198;
  wire [0:0] R1197;
  wire [0:0] R1196;
  wire [0:0] R1195;
  wire [0:0] R1194;
  wire [0:0] R1193;
  wire [0:0] R1192;
  wire [0:0] R1191;
  wire [0:0] R1190;
  wire [0:0] R1189;
  wire [0:0] R1188;
  wire [0:0] R1187;
  wire [0:0] R1186;
  wire [0:0] R1185;
  wire [0:0] R1184;
  wire [0:0] R1183;
  wire [0:0] R1182;
  wire [0:0] R1181;
  wire [0:0] R1180;
  wire [0:0] R1179;
  wire [0:0] R1178;
  wire [0:0] R1177;
  wire [0:0] R1176;
  wire [0:0] R1175;
  wire [0:0] R1174;
  wire [0:0] R1173;
  wire [0:0] R1172;
  wire [0:0] R1171;
  wire [0:0] R1170;
  wire [0:0] R1169;
  wire [0:0] R1168;
  wire [0:0] R1167;
  wire [0:0] R1166;
  wire [0:0] R1165;
  wire [0:0] R1164;
  wire [0:0] R1163;
  wire [0:0] R1162;
  wire [0:0] R1161;
  wire [0:0] R1160;
  wire [0:0] R1159;
  wire [0:0] R1158;
  wire [0:0] R1157;
  wire [0:0] R1156;
  wire [0:0] R1155;
  wire [0:0] R1154;
  wire [0:0] R1153;
  wire [0:0] R1152;
  wire [0:0] R1151;
  wire [0:0] R1150;
  wire [0:0] R1149;
  wire [0:0] R1148;
  wire [0:0] R1147;
  wire [0:0] R1146;
  wire [0:0] R1145;
  wire [0:0] R1144;
  wire [0:0] R1143;
  wire [0:0] R1142;
  wire [0:0] R1141;
  wire [0:0] R1140;
  wire [0:0] R1139;
  wire [0:0] R1138;
  wire [0:0] R1137;
  wire [0:0] R1136;
  wire [0:0] R1135;
  wire [0:0] R1134;
  wire [0:0] R1133;
  wire [0:0] R1132;
  wire [0:0] R1131;
  wire [0:0] R1130;
  wire [0:0] R1129;
  wire [0:0] R1128;
  wire [0:0] R1127;
  wire [0:0] R1126;
  wire [0:0] R1125;
  wire [0:0] R1124;
  wire [0:0] R1123;
  wire [0:0] R1122;
  wire [31:0] R1121;
  wire [63:0] R1120;
  wire [63:0] R1119;
  wire [31:0] R1118;
  wire [31:0] R1117;
  wire [31:0] R1116;
  wire [31:0] R1115;
  wire [31:0] R1114;
  wire [31:0] R1113;
  wire [31:0] R1112;
  wire [31:0] R1111;
  wire [31:0] R1110;
  wire [31:0] R1109;
  wire [31:0] R1108;
  wire [31:0] R1107;
  wire [31:0] R1106;
  wire [31:0] R1105;
  wire [31:0] R1104;
  wire [31:0] R1103;
  wire [31:0] R1102;
  wire [31:0] R1101;
  wire [31:0] R1100;
  wire [31:0] R1099;
  wire [31:0] R1098;
  wire [31:0] R1097;
  wire [31:0] R1096;
  wire [31:0] R1095;
  wire [31:0] R1094;
  wire [31:0] R1093;
  wire [31:0] R1092;
  wire [31:0] R1091;
  wire [31:0] R1090;
  wire [31:0] R1089;
  wire [31:0] R1088;
  wire [31:0] R1087;
  wire [31:0] R1086;
  wire [31:0] R1085;
  wire [31:0] R1084;
  wire [31:0] R1083;
  wire [31:0] R1082;
  wire [31:0] R1081;
  wire [31:0] R1080;
  wire [31:0] R1079;
  wire [31:0] R1078;
  wire [31:0] R1077;
  wire [31:0] R1076;
  wire [31:0] R1075;
  wire [31:0] R1074;
  wire [31:0] R1073;
  wire [31:0] R1072;
  wire [31:0] R1071;
  wire [31:0] R1070;
  wire [31:0] R1069;
  wire [31:0] R1068;
  wire [31:0] R1067;
  wire [31:0] R1066;
  wire [31:0] R1065;
  wire [31:0] R1064;
  wire [31:0] R1063;
  wire [31:0] R1062;
  wire [31:0] R1061;
  wire [31:0] R1060;
  wire [31:0] R1059;
  wire [31:0] R1058;
  wire [31:0] R1057;
  wire [31:0] R1056;
  wire [31:0] R1055;
  wire [31:0] R1054;
  wire [31:0] R1053;
  wire [31:0] R1052;
  wire [31:0] R1051;
  wire [31:0] R1050;
  wire [31:0] R1049;
  wire [31:0] R1048;
  wire [31:0] R1047;
  wire [31:0] R1046;
  wire [31:0] R1045;
  wire [31:0] R1044;
  wire [31:0] R1043;
  wire [31:0] R1042;
  wire [31:0] R1041;
  wire [31:0] R1040;
  wire [31:0] R1039;
  wire [31:0] R1038;
  wire [31:0] R1037;
  wire [31:0] R1036;
  wire [31:0] R1035;
  wire [31:0] R1034;
  wire [31:0] R1033;
  wire [31:0] R1032;
  wire [31:0] R1031;
  wire [31:0] R1030;
  wire [31:0] R1029;
  wire [31:0] R1028;
  wire [31:0] R1027;
  wire [31:0] R1026;
  wire [31:0] R1025;
  wire [31:0] R1024;
  wire [31:0] R1023;
  wire [31:0] R1022;
  wire [31:0] R1021;
  wire [31:0] R1020;
  wire [31:0] R1019;
  wire [31:0] R1018;
  wire [31:0] R1017;
  wire [31:0] R1016;
  wire [31:0] R1015;
  wire [63:0] R1014;
  wire [63:0] R1013;
  wire [0:0] R1012;
  wire [0:0] R1011;
  wire [0:0] R1010;
  wire [0:0] R1009;
  wire [0:0] R1008;
  wire [0:0] R1007;
  wire [0:0] R1006;
  wire [0:0] R1005;
  wire [0:0] R1004;
  wire [0:0] R1003;
  wire [0:0] R1002;
  wire [0:0] R1001;
  wire [0:0] R1000;
  wire [0:0] R999;
  wire [0:0] R998;
  wire [0:0] R997;
  wire [0:0] R996;
  wire [0:0] R995;
  wire [0:0] R994;
  wire [0:0] R993;
  wire [0:0] R992;
  wire [0:0] R991;
  wire [0:0] R990;
  wire [0:0] R989;
  wire [0:0] R988;
  wire [0:0] R987;
  wire [0:0] R986;
  wire [0:0] R985;
  wire [0:0] R984;
  wire [0:0] R983;
  wire [0:0] R982;
  wire [0:0] R981;
  wire [0:0] R980;
  wire [0:0] R979;
  wire [0:0] R978;
  wire [0:0] R977;
  wire [0:0] R976;
  wire [0:0] R975;
  wire [0:0] R974;
  wire [0:0] R973;
  wire [0:0] R972;
  wire [0:0] R971;
  wire [0:0] R970;
  wire [0:0] R969;
  wire [0:0] R968;
  wire [0:0] R967;
  wire [0:0] R966;
  wire [0:0] R965;
  wire [0:0] R964;
  wire [0:0] R963;
  wire [0:0] R962;
  wire [0:0] R961;
  wire [0:0] R960;
  wire [0:0] R959;
  wire [0:0] R958;
  wire [0:0] R957;
  wire [0:0] R956;
  wire [0:0] R955;
  wire [0:0] R954;
  wire [0:0] R953;
  wire [0:0] R952;
  wire [0:0] R951;
  wire [0:0] R950;
  wire [0:0] R949;
  wire [0:0] R948;
  wire [0:0] R947;
  wire [0:0] R946;
  wire [0:0] R945;
  wire [0:0] R944;
  wire [0:0] R943;
  wire [0:0] R942;
  wire [0:0] R941;
  wire [0:0] R940;
  wire [0:0] R939;
  wire [0:0] R938;
  wire [0:0] R937;
  wire [0:0] R936;
  wire [0:0] R935;
  wire [0:0] R934;
  wire [0:0] R933;
  wire [0:0] R932;
  wire [0:0] R931;
  wire [0:0] R930;
  wire [0:0] R929;
  wire [0:0] R928;
  wire [0:0] R927;
  wire [0:0] R926;
  wire [0:0] R925;
  wire [0:0] R924;
  wire [0:0] R923;
  wire [0:0] R922;
  wire [0:0] R921;
  wire [0:0] R920;
  wire [0:0] R919;
  wire [0:0] R918;
  wire [0:0] R917;
  wire [0:0] R916;
  wire [0:0] R915;
  wire [0:0] R914;
  wire [0:0] R913;
  wire [0:0] R912;
  wire [0:0] R911;
  wire [0:0] R910;
  wire [0:0] R909;
  wire [0:0] R908;
  wire [0:0] R907;
  wire [0:0] R906;
  wire [0:0] R905;
  wire [31:0] R904;
  wire [63:0] R903;
  wire [63:0] R902;
  wire [31:0] R901;
  wire [31:0] R900;
  wire [31:0] R899;
  wire [31:0] R898;
  wire [31:0] R897;
  wire [31:0] R896;
  wire [31:0] R895;
  wire [31:0] R894;
  wire [31:0] R893;
  wire [31:0] R892;
  wire [31:0] R891;
  wire [31:0] R890;
  wire [31:0] R889;
  wire [31:0] R888;
  wire [31:0] R887;
  wire [31:0] R886;
  wire [31:0] R885;
  wire [31:0] R884;
  wire [31:0] R883;
  wire [31:0] R882;
  wire [31:0] R881;
  wire [31:0] R880;
  wire [31:0] R879;
  wire [31:0] R878;
  wire [31:0] R877;
  wire [31:0] R876;
  wire [31:0] R875;
  wire [31:0] R874;
  wire [31:0] R873;
  wire [31:0] R872;
  wire [31:0] R871;
  wire [31:0] R870;
  wire [31:0] R869;
  wire [31:0] R868;
  wire [31:0] R867;
  wire [31:0] R866;
  wire [31:0] R865;
  wire [31:0] R864;
  wire [31:0] R863;
  wire [31:0] R862;
  wire [31:0] R861;
  wire [31:0] R860;
  wire [31:0] R859;
  wire [31:0] R858;
  wire [31:0] R857;
  wire [31:0] R856;
  wire [31:0] R855;
  wire [31:0] R854;
  wire [31:0] R853;
  wire [31:0] R852;
  wire [31:0] R851;
  wire [31:0] R850;
  wire [31:0] R849;
  wire [31:0] R848;
  wire [31:0] R847;
  wire [31:0] R846;
  wire [31:0] R845;
  wire [31:0] R844;
  wire [31:0] R843;
  wire [31:0] R842;
  wire [31:0] R841;
  wire [31:0] R840;
  wire [31:0] R839;
  wire [31:0] R838;
  wire [31:0] R837;
  wire [31:0] R836;
  wire [31:0] R835;
  wire [31:0] R834;
  wire [31:0] R833;
  wire [31:0] R832;
  wire [31:0] R831;
  wire [31:0] R830;
  wire [31:0] R829;
  wire [31:0] R828;
  wire [31:0] R827;
  wire [31:0] R826;
  wire [31:0] R825;
  wire [31:0] R824;
  wire [31:0] R823;
  wire [31:0] R822;
  wire [31:0] R821;
  wire [31:0] R820;
  wire [31:0] R819;
  wire [31:0] R818;
  wire [31:0] R817;
  wire [31:0] R816;
  wire [31:0] R815;
  wire [31:0] R814;
  wire [31:0] R813;
  wire [31:0] R812;
  wire [31:0] R811;
  wire [31:0] R810;
  wire [31:0] R809;
  wire [31:0] R808;
  wire [31:0] R807;
  wire [31:0] R806;
  wire [31:0] R805;
  wire [31:0] R804;
  wire [31:0] R803;
  wire [31:0] R802;
  wire [31:0] R801;
  wire [31:0] R800;
  wire [31:0] R799;
  wire [31:0] R798;
  wire [31:0] R797;
  wire [31:0] R796;
  wire [31:0] R795;
  wire [31:0] R794;
  wire [31:0] R793;
  wire [31:0] R792;
  wire [31:0] R791;
  wire [31:0] R790;
  wire [31:0] R789;
  wire [63:0] R788;
  wire [63:0] R787;
  wire [0:0] R786;
  wire [0:0] R785;
  wire [0:0] R784;
  wire [0:0] R783;
  wire [0:0] R782;
  wire [0:0] R781;
  wire [0:0] R780;
  wire [0:0] R779;
  wire [0:0] R778;
  wire [0:0] R777;
  wire [0:0] R776;
  wire [0:0] R775;
  wire [0:0] R774;
  wire [0:0] R773;
  wire [0:0] R772;
  wire [0:0] R771;
  wire [0:0] R770;
  wire [0:0] R769;
  wire [0:0] R768;
  wire [0:0] R767;
  wire [0:0] R766;
  wire [0:0] R765;
  wire [0:0] R764;
  wire [0:0] R763;
  wire [0:0] R762;
  wire [0:0] R761;
  wire [0:0] R760;
  wire [0:0] R759;
  wire [0:0] R758;
  wire [0:0] R757;
  wire [0:0] R756;
  wire [0:0] R755;
  wire [0:0] R754;
  wire [0:0] R753;
  wire [0:0] R752;
  wire [0:0] R751;
  wire [0:0] R750;
  wire [0:0] R749;
  wire [0:0] R748;
  wire [0:0] R747;
  wire [0:0] R746;
  wire [0:0] R745;
  wire [0:0] R744;
  wire [0:0] R743;
  wire [0:0] R742;
  wire [0:0] R741;
  wire [0:0] R740;
  wire [0:0] R739;
  wire [0:0] R738;
  wire [0:0] R737;
  wire [0:0] R736;
  wire [0:0] R735;
  wire [0:0] R734;
  wire [0:0] R733;
  wire [0:0] R732;
  wire [0:0] R731;
  wire [0:0] R730;
  wire [0:0] R729;
  wire [0:0] R728;
  wire [0:0] R727;
  wire [0:0] R726;
  wire [0:0] R725;
  wire [0:0] R724;
  wire [0:0] R723;
  wire [0:0] R722;
  wire [0:0] R721;
  wire [0:0] R720;
  wire [0:0] R719;
  wire [0:0] R718;
  wire [0:0] R717;
  wire [0:0] R716;
  wire [0:0] R715;
  wire [0:0] R714;
  wire [0:0] R713;
  wire [0:0] R712;
  wire [0:0] R711;
  wire [0:0] R710;
  wire [0:0] R709;
  wire [0:0] R708;
  wire [0:0] R707;
  wire [0:0] R706;
  wire [0:0] R705;
  wire [0:0] R704;
  wire [0:0] R703;
  wire [0:0] R702;
  wire [0:0] R701;
  wire [0:0] R700;
  wire [0:0] R699;
  wire [0:0] R698;
  wire [0:0] R697;
  wire [0:0] R696;
  wire [0:0] R695;
  wire [0:0] R694;
  wire [0:0] R693;
  wire [0:0] R692;
  wire [0:0] R691;
  wire [0:0] R690;
  wire [0:0] R689;
  wire [0:0] R688;
  wire [0:0] R687;
  wire [0:0] R686;
  wire [0:0] R685;
  wire [0:0] R684;
  wire [0:0] R683;
  wire [0:0] R682;
  wire [0:0] R681;
  wire [0:0] R680;
  wire [0:0] R679;
  wire [0:0] R678;
  wire [0:0] R677;
  wire [0:0] R676;
  wire [0:0] R675;
  wire [0:0] R674;
  wire [0:0] R673;
  wire [0:0] R672;
  wire [0:0] R671;
  wire [0:0] R670;
  wire [31:0] R669;
  wire [63:0] R668;
  wire [63:0] R667;
  wire [31:0] R666;
  wire [31:0] R665;
  wire [31:0] R664;
  wire [31:0] R663;
  wire [31:0] R662;
  wire [31:0] R661;
  wire [31:0] R660;
  wire [31:0] R659;
  wire [31:0] R658;
  wire [31:0] R657;
  wire [31:0] R656;
  wire [31:0] R655;
  wire [31:0] R654;
  wire [31:0] R653;
  wire [31:0] R652;
  wire [31:0] R651;
  wire [31:0] R650;
  wire [31:0] R649;
  wire [31:0] R648;
  wire [31:0] R647;
  wire [31:0] R646;
  wire [31:0] R645;
  wire [31:0] R644;
  wire [31:0] R643;
  wire [31:0] R642;
  wire [31:0] R641;
  wire [31:0] R640;
  wire [31:0] R639;
  wire [31:0] R638;
  wire [31:0] R637;
  wire [31:0] R636;
  wire [31:0] R635;
  wire [31:0] R634;
  wire [31:0] R633;
  wire [31:0] R632;
  wire [31:0] R631;
  wire [31:0] R630;
  wire [31:0] R629;
  wire [31:0] R628;
  wire [31:0] R627;
  wire [31:0] R626;
  wire [31:0] R625;
  wire [31:0] R624;
  wire [31:0] R623;
  wire [31:0] R622;
  wire [31:0] R621;
  wire [31:0] R620;
  wire [31:0] R619;
  wire [31:0] R618;
  wire [31:0] R617;
  wire [31:0] R616;
  wire [31:0] R615;
  wire [31:0] R614;
  wire [31:0] R613;
  wire [31:0] R612;
  wire [31:0] R611;
  wire [31:0] R610;
  wire [31:0] R609;
  wire [31:0] R608;
  wire [31:0] R607;
  wire [31:0] R606;
  wire [31:0] R605;
  wire [31:0] R604;
  wire [31:0] R603;
  wire [31:0] R602;
  wire [31:0] R601;
  wire [31:0] R600;
  wire [31:0] R599;
  wire [31:0] R598;
  wire [31:0] R597;
  wire [31:0] R596;
  wire [31:0] R595;
  wire [31:0] R594;
  wire [31:0] R593;
  wire [31:0] R592;
  wire [31:0] R591;
  wire [31:0] R590;
  wire [31:0] R589;
  wire [31:0] R588;
  wire [31:0] R587;
  wire [31:0] R586;
  wire [31:0] R585;
  wire [31:0] R584;
  wire [31:0] R583;
  wire [31:0] R582;
  wire [31:0] R581;
  wire [31:0] R580;
  wire [31:0] R579;
  wire [31:0] R578;
  wire [31:0] R577;
  wire [31:0] R576;
  wire [31:0] R575;
  wire [31:0] R574;
  wire [31:0] R573;
  wire [31:0] R572;
  wire [31:0] R571;
  wire [31:0] R570;
  wire [31:0] R569;
  wire [31:0] R568;
  wire [31:0] R567;
  wire [31:0] R566;
  wire [31:0] R565;
  wire [31:0] R564;
  wire [31:0] R563;
  wire [31:0] R562;
  wire [31:0] R561;
  wire [31:0] R560;
  wire [31:0] R559;
  wire [31:0] R558;
  wire [31:0] R557;
  wire [31:0] R556;
  wire [31:0] R555;
  wire [31:0] R554;
  wire [31:0] R553;
  wire [31:0] R552;
  wire [31:0] R551;
  wire [31:0] R550;
  wire [31:0] R549;
  wire [31:0] R548;
  wire [31:0] R547;
  wire [31:0] R546;
  wire [15:0] R545;
  wire [63:0] R544;
  wire [63:0] R543;
  wire [0:0] R542;
  wire [0:0] R541;
  wire [0:0] R540;
  wire [0:0] R539;
  wire [0:0] R538;
  wire [0:0] R537;
  wire [0:0] R536;
  wire [0:0] R535;
  wire [0:0] R534;
  wire [0:0] R533;
  wire [0:0] R532;
  wire [0:0] R531;
  wire [0:0] R530;
  wire [0:0] R529;
  wire [0:0] R528;
  wire [0:0] R527;
  wire [0:0] R526;
  wire [0:0] R525;
  wire [0:0] R524;
  wire [0:0] R523;
  wire [0:0] R522;
  wire [0:0] R521;
  wire [0:0] R520;
  wire [0:0] R519;
  wire [0:0] R518;
  wire [0:0] R517;
  wire [0:0] R516;
  wire [0:0] R515;
  wire [0:0] R514;
  wire [0:0] R513;
  wire [0:0] R512;
  wire [0:0] R511;
  wire [0:0] R510;
  wire [0:0] R509;
  wire [0:0] R508;
  wire [0:0] R507;
  wire [0:0] R506;
  wire [0:0] R505;
  wire [0:0] R504;
  wire [0:0] R503;
  wire [0:0] R502;
  wire [0:0] R501;
  wire [0:0] R500;
  wire [0:0] R499;
  wire [0:0] R498;
  wire [0:0] R497;
  wire [0:0] R496;
  wire [0:0] R495;
  wire [0:0] R494;
  wire [0:0] R493;
  wire [0:0] R492;
  wire [0:0] R491;
  wire [0:0] R490;
  wire [0:0] R489;
  wire [0:0] R488;
  wire [0:0] R487;
  wire [0:0] R486;
  wire [0:0] R485;
  wire [0:0] R484;
  wire [0:0] R483;
  wire [0:0] R482;
  wire [0:0] R481;
  wire [0:0] R480;
  wire [0:0] R479;
  wire [0:0] R478;
  wire [0:0] R477;
  wire [0:0] R476;
  wire [0:0] R475;
  wire [0:0] R474;
  wire [0:0] R473;
  wire [0:0] R472;
  wire [0:0] R471;
  wire [0:0] R470;
  wire [0:0] R469;
  wire [0:0] R468;
  wire [0:0] R467;
  wire [0:0] R466;
  wire [0:0] R465;
  wire [0:0] R464;
  wire [0:0] R463;
  wire [0:0] R462;
  wire [0:0] R461;
  wire [0:0] R460;
  wire [0:0] R459;
  wire [0:0] R458;
  wire [0:0] R457;
  wire [0:0] R456;
  wire [0:0] R455;
  wire [0:0] R454;
  wire [0:0] R453;
  wire [0:0] R452;
  wire [0:0] R451;
  wire [0:0] R450;
  wire [0:0] R449;
  wire [0:0] R448;
  wire [0:0] R447;
  wire [0:0] R446;
  wire [0:0] R445;
  wire [0:0] R444;
  wire [0:0] R443;
  wire [0:0] R442;
  wire [0:0] R441;
  wire [0:0] R440;
  wire [0:0] R439;
  wire [0:0] R438;
  wire [0:0] R437;
  wire [0:0] R436;
  wire [0:0] R435;
  wire [0:0] R434;
  wire [0:0] R433;
  wire [0:0] R432;
  wire [0:0] R431;
  wire [0:0] R430;
  wire [0:0] R429;
  wire [0:0] R428;
  wire [0:0] R427;
  wire [0:0] R426;
  wire [0:0] R425;
  wire [0:0] R424;
  wire [0:0] R423;
  wire [0:0] R422;
  wire [0:0] R421;
  wire [0:0] R420;
  wire [0:0] R419;
  wire [0:0] R418;
  wire [0:0] R417;
  wire [15:0] R416;
  wire [63:0] R415;
  wire [63:0] R414;
  wire [31:0] R413;
  wire [31:0] R412;
  wire [31:0] R411;
  wire [31:0] R410;
  wire [31:0] R409;
  wire [31:0] R408;
  wire [31:0] R407;
  wire [31:0] R406;
  wire [31:0] R405;
  wire [31:0] R404;
  wire [31:0] R403;
  wire [31:0] R402;
  wire [31:0] R401;
  wire [31:0] R400;
  wire [31:0] R399;
  wire [31:0] R398;
  wire [31:0] R397;
  wire [31:0] R396;
  wire [31:0] R395;
  wire [31:0] R394;
  wire [31:0] R393;
  wire [31:0] R392;
  wire [31:0] R391;
  wire [31:0] R390;
  wire [31:0] R389;
  wire [31:0] R388;
  wire [31:0] R387;
  wire [31:0] R386;
  wire [31:0] R385;
  wire [31:0] R384;
  wire [31:0] R383;
  wire [31:0] R382;
  wire [31:0] R381;
  wire [31:0] R380;
  wire [31:0] R379;
  wire [31:0] R378;
  wire [31:0] R377;
  wire [31:0] R376;
  wire [31:0] R375;
  wire [31:0] R374;
  wire [31:0] R373;
  wire [31:0] R372;
  wire [31:0] R371;
  wire [31:0] R370;
  wire [31:0] R369;
  wire [31:0] R368;
  wire [31:0] R367;
  wire [31:0] R366;
  wire [31:0] R365;
  wire [31:0] R364;
  wire [31:0] R363;
  wire [31:0] R362;
  wire [31:0] R361;
  wire [31:0] R360;
  wire [31:0] R359;
  wire [31:0] R358;
  wire [31:0] R357;
  wire [31:0] R356;
  wire [31:0] R355;
  wire [31:0] R354;
  wire [31:0] R353;
  wire [31:0] R352;
  wire [31:0] R351;
  wire [31:0] R350;
  wire [31:0] R349;
  wire [31:0] R348;
  wire [31:0] R347;
  wire [31:0] R346;
  wire [31:0] R345;
  wire [31:0] R344;
  wire [31:0] R343;
  wire [31:0] R342;
  wire [31:0] R341;
  wire [31:0] R340;
  wire [31:0] R339;
  wire [31:0] R338;
  wire [31:0] R337;
  wire [31:0] R336;
  wire [31:0] R335;
  wire [31:0] R334;
  wire [31:0] R333;
  wire [31:0] R332;
  wire [31:0] R331;
  wire [31:0] R330;
  wire [31:0] R329;
  wire [31:0] R328;
  wire [31:0] R327;
  wire [31:0] R326;
  wire [31:0] R325;
  wire [31:0] R324;
  wire [31:0] R323;
  wire [31:0] R322;
  wire [31:0] R321;
  wire [31:0] R320;
  wire [31:0] R319;
  wire [31:0] R318;
  wire [31:0] R317;
  wire [31:0] R316;
  wire [31:0] R315;
  wire [31:0] R314;
  wire [31:0] R313;
  wire [31:0] R312;
  wire [31:0] R311;
  wire [31:0] R310;
  wire [31:0] R309;
  wire [31:0] R308;
  wire [31:0] R307;
  wire [31:0] R306;
  wire [31:0] R305;
  wire [31:0] R304;
  wire [31:0] R303;
  wire [31:0] R302;
  wire [31:0] R301;
  wire [31:0] R300;
  wire [31:0] R299;
  wire [31:0] R298;
  wire [31:0] R297;
  wire [31:0] R296;
  wire [31:0] R295;
  wire [31:0] R294;
  wire [31:0] R293;
  wire [31:0] R292;
  wire [31:0] R291;
  wire [31:0] R290;
  wire [31:0] R289;
  wire [31:0] R288;
  wire [31:0] R287;
  wire [31:0] R286;
  wire [7:0] mux13;
  wire [7:0] mux12;
  wire [7:0] mux11;
  wire [7:0] mux10;
  wire [7:0] mux9;
  wire [7:0] mux8;
  wire [7:0] mux7;
  wire [7:0] mux6;
  wire [7:0] mux5;
  wire [7:0] mux4;
  wire [7:0] mux3;
  wire [7:0] mux2;
  wire [7:0] mux1;
  wire [7:0] mux0;
  wire [7:0] _234;
  wire [7:0] _227;
  wire [63:0] _226;
  wire [63:0] _225;
  wire [7:0] _238;
  wire [7:0] _224;
  wire [63:0] _223;
  wire [63:0] _222;
  wire [7:0] _242;
  wire [7:0] _221;
  wire [63:0] _220;
  wire [63:0] _219;
  wire [7:0] _246;
  wire [7:0] _218;
  wire [63:0] _217;
  wire [63:0] _216;
  wire [7:0] _250;
  wire [7:0] _215;
  wire [63:0] _214;
  wire [63:0] _213;
  wire [7:0] _254;
  wire [7:0] _212;
  wire [63:0] _211;
  wire [63:0] _210;
  wire [7:0] _258;
  wire [7:0] _209;
  wire [63:0] _208;
  wire [63:0] _207;
  wire [7:0] _263;
  wire [7:0] _206;
  wire [63:0] _205;
  wire [63:0] _204;
  wire [7:0] _267;
  wire [7:0] _203;
  wire [63:0] _202;
  wire [63:0] _201;
  wire [7:0] _271;
  wire [7:0] _200;
  wire [63:0] _199;
  wire [63:0] _198;
  wire [7:0] _275;
  wire [7:0] _197;
  wire [63:0] _196;
  wire [63:0] _195;
  wire [7:0] _279;
  wire [7:0] _194;
  wire [63:0] _193;
  wire [63:0] _192;
  wire [7:0] _283;
  wire [7:0] _191;
  wire [63:0] _190;
  wire [63:0] _189;
  wire [7:0] _287;
  wire [7:0] _188;
  wire [63:0] _187;
  wire [63:0] _186;
  wire [7:0] _290;
  wire [7:0] _185;
  wire [63:0] _184;
  wire [63:0] _183;
  wire [31:0] idx_288;
  wire [31:0] _182;
  wire [31:0] _181;
  wire [31:0] _180;
  wire [31:0] _179;
  wire [31:0] _178;
  wire [63:0] _177;
  wire [63:0] _176;
  wire [63:0] _175;
  wire [0:0] ifout201;
  wire [31:0] _174;
  wire [63:0] _173;
  wire [63:0] _172;
  wire [63:0] _171;
  wire [31:0] idx_284;
  wire [31:0] _170;
  wire [31:0] _169;
  wire [63:0] _168;
  wire [31:0] _167;
  wire [31:0] _166;
  wire [31:0] _165;
  wire [63:0] _164;
  wire [63:0] _163;
  wire [63:0] _162;
  wire [0:0] ifout186;
  wire [31:0] _161;
  wire [63:0] _160;
  wire [63:0] _159;
  wire [63:0] _158;
  wire [31:0] idx_280;
  wire [31:0] _157;
  wire [31:0] _156;
  wire [63:0] _155;
  wire [31:0] _154;
  wire [31:0] _153;
  wire [31:0] _152;
  wire [63:0] _151;
  wire [63:0] _150;
  wire [63:0] _149;
  wire [0:0] ifout171;
  wire [31:0] _148;
  wire [63:0] _147;
  wire [63:0] _146;
  wire [63:0] _145;
  wire [31:0] idx_276;
  wire [31:0] _144;
  wire [31:0] _143;
  wire [63:0] _142;
  wire [31:0] _141;
  wire [31:0] _140;
  wire [31:0] _139;
  wire [63:0] _138;
  wire [63:0] _137;
  wire [63:0] _136;
  wire [0:0] ifout156;
  wire [31:0] _135;
  wire [63:0] _134;
  wire [63:0] _133;
  wire [63:0] _132;
  wire [31:0] idx_272;
  wire [31:0] _131;
  wire [31:0] _130;
  wire [63:0] _129;
  wire [31:0] _128;
  wire [31:0] _127;
  wire [31:0] _126;
  wire [63:0] _125;
  wire [63:0] _124;
  wire [63:0] _123;
  wire [0:0] ifout141;
  wire [31:0] _122;
  wire [63:0] _121;
  wire [63:0] _120;
  wire [63:0] _119;
  wire [31:0] idx_268;
  wire [31:0] _118;
  wire [31:0] _117;
  wire [63:0] _116;
  wire [31:0] _115;
  wire [31:0] _114;
  wire [31:0] _113;
  wire [63:0] _112;
  wire [63:0] _111;
  wire [63:0] _110;
  wire [0:0] ifout126;
  wire [31:0] _109;
  wire [63:0] _108;
  wire [63:0] _107;
  wire [63:0] _106;
  wire [31:0] idx_264;
  wire [31:0] _105;
  wire [31:0] _104;
  wire [63:0] _103;
  wire [31:0] _102;
  wire [31:0] _101;
  wire [31:0] _100;
  wire [63:0] _99;
  wire [63:0] _98;
  wire [63:0] _97;
  wire [0:0] ifout111;
  wire [31:0] _96;
  wire [63:0] _95;
  wire [63:0] _94;
  wire [63:0] _93;
  wire [31:0] idx_260;
  wire [31:0] _92;
  wire [63:0] _91;
  wire [31:0] _90;
  wire [31:0] _89;
  wire [31:0] _88;
  wire [63:0] _87;
  wire [63:0] _86;
  wire [63:0] _85;
  wire [0:0] ifout97;
  wire [31:0] _84;
  wire [63:0] _83;
  wire [63:0] _82;
  wire [63:0] _81;
  wire [31:0] idx_255;
  wire [31:0] _80;
  wire [31:0] _79;
  wire [31:0] _78;
  wire [31:0] _77;
  wire [31:0] _76;
  wire [63:0] _75;
  wire [63:0] _74;
  wire [63:0] _73;
  wire [0:0] ifout83;
  wire [31:0] _72;
  wire [63:0] _71;
  wire [63:0] _70;
  wire [63:0] _69;
  wire [31:0] idx_251;
  wire [31:0] _68;
  wire [31:0] _67;
  wire [63:0] _66;
  wire [31:0] _65;
  wire [31:0] _64;
  wire [31:0] _63;
  wire [63:0] _62;
  wire [63:0] _61;
  wire [63:0] _60;
  wire [0:0] ifout68;
  wire [31:0] _59;
  wire [63:0] _58;
  wire [63:0] _57;
  wire [63:0] _56;
  wire [31:0] idx_247;
  wire [31:0] _55;
  wire [31:0] _54;
  wire [63:0] _53;
  wire [31:0] _52;
  wire [31:0] _51;
  wire [31:0] _50;
  wire [63:0] _49;
  wire [63:0] _48;
  wire [63:0] _47;
  wire [0:0] ifout53;
  wire [31:0] _46;
  wire [63:0] _45;
  wire [63:0] _44;
  wire [63:0] _43;
  wire [31:0] idx_243;
  wire [31:0] _42;
  wire [31:0] _41;
  wire [63:0] _40;
  wire [31:0] _39;
  wire [31:0] _38;
  wire [31:0] _37;
  wire [63:0] _36;
  wire [63:0] _35;
  wire [63:0] _34;
  wire [0:0] ifout38;
  wire [31:0] _33;
  wire [63:0] _32;
  wire [63:0] _31;
  wire [63:0] _30;
  wire [31:0] idx_239;
  wire [31:0] _29;
  wire [31:0] _28;
  wire [63:0] _27;
  wire [31:0] _26;
  wire [31:0] _25;
  wire [31:0] _24;
  wire [63:0] _23;
  wire [63:0] _22;
  wire [63:0] _21;
  wire [0:0] ifout23;
  wire [31:0] _20;
  wire [63:0] _19;
  wire [63:0] _18;
  wire [63:0] _17;
  wire [31:0] idx_235;
  wire [31:0] _16;
  wire [31:0] _15;
  wire [63:0] _14;
  wire [31:0] _13;
  wire [31:0] _12;
  wire [31:0] _11;
  wire [31:0] _10;
  wire [15:0] _9;
  wire [63:0] _8;
  wire [63:0] _7;
  wire [63:0] _6;
  wire [0:0] ifout6;
  wire [15:0] _5;
  wire [63:0] _4;
  wire [63:0] _3;
  wire [63:0] _2;
  wire [31:0] idx_230;
  wire [63:0] _1;
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op0 (.out1(_1), .in1(ip1_229_D), .in2(6 'd 48));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1 (.out1(idx_230), .in1(_1));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op285 (.out1(R286), .clock(clock), .in1(idx_230));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2 (.out1(_2), .in1(R286));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op3 (.out1(_3), .in1(_2), .in2(1 'd 1));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op286 (.out1(R287), .clock(clock), .in1(R286));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op413 (.out1(R414), .clock(clock), .in1(_3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op4 (.out1(_4), .in1(C16_231_D), .in2(R414));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op287 (.out1(R288), .clock(clock), .in1(R287));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op414 (.out1(R415), .clock(clock), .in1(_4));
  SRAM op5 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_5),.ADR(R415));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op288 (.out1(R289), .clock(clock), .in1(R288));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op415 (.out1(R416), .clock(clock), .in1(_5));
  NE_EXPR #(.BITSIZE_in1(16), .BITSIZE_in2(1),.BITSIZE_out1(1)) op6 (.out1(ifout6), .in1(R416), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op7 (.out1(_6), .in1(R289));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op8 (.out1(_7), .in1(_6), .in2(1 'd 1));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op289 (.out1(R290), .clock(clock), .in1(R289));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op416 (.out1(R417), .clock(clock), .in1(ifout6));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op542 (.out1(R543), .clock(clock), .in1(_7));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op9 (.out1(_8), .in1(C16_231_D), .in2(R543));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op290 (.out1(R291), .clock(clock), .in1(R290));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op417 (.out1(R418), .clock(clock), .in1(R417));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op543 (.out1(R544), .clock(clock), .in1(_8));
  SRAM op10 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_9),.ADR(R544));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op291 (.out1(R292), .clock(clock), .in1(R291));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op418 (.out1(R419), .clock(clock), .in1(R418));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op544 (.out1(R545), .clock(clock), .in1(_9));
  cast #(.BITSIZE_in1(16), .BITSIZE_out1(32)) op11 (.out1(_10), .in1(R545));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(1), .BITSIZE_out1(32)) op12 (.out1(_11), .in1(_10), .in2(-1 'd 1));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op292 (.out1(R293), .clock(clock), .in1(R292));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op419 (.out1(R420), .clock(clock), .in1(R419));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op545 (.out1(R546), .clock(clock), .in1(_11));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(4), .BITSIZE_out1(32), .PRECISION(32)) op13 (.out1(_12), .in1(R546), .in2(4 'd 8));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op293 (.out1(R294), .clock(clock), .in1(R293));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op420 (.out1(R421), .clock(clock), .in1(R420));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op546 (.out1(R547), .clock(clock), .in1(_12));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op15 (.out1(_14), .in1(ip1_229_D), .in2(6 'd 40));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op16 (.out1(_15), .in1(_14));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op14 (.out1(_13), .in1(R547));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(8), .BITSIZE_out1(32)) op17 (.out1(_16), .in1(_15), .in2(8 'd 255));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op18 (.out1(idx_235), .in1(_13), .in2(_16));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op294 (.out1(R295), .clock(clock), .in1(R294));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op421 (.out1(R422), .clock(clock), .in1(R421));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op547 (.out1(R548), .clock(clock), .in1(idx_235));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op19 (.out1(_17), .in1(R548));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op20 (.out1(_18), .in1(_17), .in2(2 'd 2));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op295 (.out1(R296), .clock(clock), .in1(R295));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op422 (.out1(R423), .clock(clock), .in1(R422));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op548 (.out1(R549), .clock(clock), .in1(R548));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op666 (.out1(R667), .clock(clock), .in1(_18));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op21 (.out1(_19), .in1(C24_236_D), .in2(R667));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op296 (.out1(R297), .clock(clock), .in1(R296));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op423 (.out1(R424), .clock(clock), .in1(R423));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op549 (.out1(R550), .clock(clock), .in1(R549));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op667 (.out1(R668), .clock(clock), .in1(_19));
  SRAM op22 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_20),.ADR(R668));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op297 (.out1(R298), .clock(clock), .in1(R297));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op424 (.out1(R425), .clock(clock), .in1(R424));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op550 (.out1(R551), .clock(clock), .in1(R550));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op668 (.out1(R669), .clock(clock), .in1(_20));
  NE_EXPR #(.BITSIZE_in1(32), .BITSIZE_in2(1),.BITSIZE_out1(1)) op23 (.out1(ifout23), .in1(R669), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op24 (.out1(_21), .in1(R551));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op25 (.out1(_22), .in1(_21), .in2(2 'd 2));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op298 (.out1(R299), .clock(clock), .in1(R298));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op425 (.out1(R426), .clock(clock), .in1(R425));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op551 (.out1(R552), .clock(clock), .in1(R551));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op669 (.out1(R670), .clock(clock), .in1(ifout23));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op786 (.out1(R787), .clock(clock), .in1(_22));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op26 (.out1(_23), .in1(C24_236_D), .in2(R787));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op299 (.out1(R300), .clock(clock), .in1(R299));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op426 (.out1(R427), .clock(clock), .in1(R426));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op552 (.out1(R553), .clock(clock), .in1(R552));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op670 (.out1(R671), .clock(clock), .in1(R670));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op787 (.out1(R788), .clock(clock), .in1(_23));
  SRAM op27 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_24),.ADR(R788));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op300 (.out1(R301), .clock(clock), .in1(R300));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op427 (.out1(R428), .clock(clock), .in1(R427));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op553 (.out1(R554), .clock(clock), .in1(R553));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op671 (.out1(R672), .clock(clock), .in1(R671));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op788 (.out1(R789), .clock(clock), .in1(_24));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op28 (.out1(_25), .in1(R789), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op301 (.out1(R302), .clock(clock), .in1(R301));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op428 (.out1(R429), .clock(clock), .in1(R428));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op554 (.out1(R555), .clock(clock), .in1(R554));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op672 (.out1(R673), .clock(clock), .in1(R672));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op789 (.out1(R790), .clock(clock), .in1(_25));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(4), .BITSIZE_out1(32), .PRECISION(32)) op29 (.out1(_26), .in1(R790), .in2(4 'd 8));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op302 (.out1(R303), .clock(clock), .in1(R302));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op429 (.out1(R430), .clock(clock), .in1(R429));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op555 (.out1(R556), .clock(clock), .in1(R555));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op673 (.out1(R674), .clock(clock), .in1(R673));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op790 (.out1(R791), .clock(clock), .in1(_26));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op30 (.out1(_27), .in1(ip1_229_D), .in2(6 'd 32));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op31 (.out1(_28), .in1(_27));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(8), .BITSIZE_out1(32)) op32 (.out1(_29), .in1(_28), .in2(8 'd 255));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op33 (.out1(idx_239), .in1(R791), .in2(_29));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op303 (.out1(R304), .clock(clock), .in1(R303));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op430 (.out1(R431), .clock(clock), .in1(R430));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op556 (.out1(R557), .clock(clock), .in1(R556));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op674 (.out1(R675), .clock(clock), .in1(R674));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op791 (.out1(R792), .clock(clock), .in1(idx_239));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op34 (.out1(_30), .in1(R792));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op35 (.out1(_31), .in1(_30), .in2(2 'd 2));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op304 (.out1(R305), .clock(clock), .in1(R304));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op431 (.out1(R432), .clock(clock), .in1(R431));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op557 (.out1(R558), .clock(clock), .in1(R557));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op675 (.out1(R676), .clock(clock), .in1(R675));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op792 (.out1(R793), .clock(clock), .in1(R792));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op901 (.out1(R902), .clock(clock), .in1(_31));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op36 (.out1(_32), .in1(C32_240_D), .in2(R902));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op305 (.out1(R306), .clock(clock), .in1(R305));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op432 (.out1(R433), .clock(clock), .in1(R432));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op558 (.out1(R559), .clock(clock), .in1(R558));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op676 (.out1(R677), .clock(clock), .in1(R676));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op793 (.out1(R794), .clock(clock), .in1(R793));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op902 (.out1(R903), .clock(clock), .in1(_32));
  SRAM op37 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_33),.ADR(R903));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op306 (.out1(R307), .clock(clock), .in1(R306));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op433 (.out1(R434), .clock(clock), .in1(R433));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op559 (.out1(R560), .clock(clock), .in1(R559));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op677 (.out1(R678), .clock(clock), .in1(R677));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op794 (.out1(R795), .clock(clock), .in1(R794));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op903 (.out1(R904), .clock(clock), .in1(_33));
  NE_EXPR #(.BITSIZE_in1(32), .BITSIZE_in2(1),.BITSIZE_out1(1)) op38 (.out1(ifout38), .in1(R904), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op39 (.out1(_34), .in1(R795));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op40 (.out1(_35), .in1(_34), .in2(2 'd 2));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op307 (.out1(R308), .clock(clock), .in1(R307));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op434 (.out1(R435), .clock(clock), .in1(R434));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op560 (.out1(R561), .clock(clock), .in1(R560));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op678 (.out1(R679), .clock(clock), .in1(R678));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op795 (.out1(R796), .clock(clock), .in1(R795));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op904 (.out1(R905), .clock(clock), .in1(ifout38));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op1012 (.out1(R1013), .clock(clock), .in1(_35));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op41 (.out1(_36), .in1(C32_240_D), .in2(R1013));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op308 (.out1(R309), .clock(clock), .in1(R308));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op435 (.out1(R436), .clock(clock), .in1(R435));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op561 (.out1(R562), .clock(clock), .in1(R561));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op679 (.out1(R680), .clock(clock), .in1(R679));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op796 (.out1(R797), .clock(clock), .in1(R796));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op905 (.out1(R906), .clock(clock), .in1(R905));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op1013 (.out1(R1014), .clock(clock), .in1(_36));
  SRAM op42 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_37),.ADR(R1014));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op309 (.out1(R310), .clock(clock), .in1(R309));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op436 (.out1(R437), .clock(clock), .in1(R436));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op562 (.out1(R563), .clock(clock), .in1(R562));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op680 (.out1(R681), .clock(clock), .in1(R680));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op797 (.out1(R798), .clock(clock), .in1(R797));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op906 (.out1(R907), .clock(clock), .in1(R906));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1014 (.out1(R1015), .clock(clock), .in1(_37));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op43 (.out1(_38), .in1(R1015), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op310 (.out1(R311), .clock(clock), .in1(R310));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op437 (.out1(R438), .clock(clock), .in1(R437));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op563 (.out1(R564), .clock(clock), .in1(R563));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op681 (.out1(R682), .clock(clock), .in1(R681));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op798 (.out1(R799), .clock(clock), .in1(R798));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op907 (.out1(R908), .clock(clock), .in1(R907));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1015 (.out1(R1016), .clock(clock), .in1(_38));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(4), .BITSIZE_out1(32), .PRECISION(32)) op44 (.out1(_39), .in1(R1016), .in2(4 'd 8));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op311 (.out1(R312), .clock(clock), .in1(R311));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op438 (.out1(R439), .clock(clock), .in1(R438));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op564 (.out1(R565), .clock(clock), .in1(R564));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op682 (.out1(R683), .clock(clock), .in1(R682));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op799 (.out1(R800), .clock(clock), .in1(R799));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op908 (.out1(R909), .clock(clock), .in1(R908));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1016 (.out1(R1017), .clock(clock), .in1(_39));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(5), .BITSIZE_out1(64), .PRECISION(64)) op45 (.out1(_40), .in1(ip1_229_D), .in2(5 'd 24));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op46 (.out1(_41), .in1(_40));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(8), .BITSIZE_out1(32)) op47 (.out1(_42), .in1(_41), .in2(8 'd 255));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op48 (.out1(idx_243), .in1(R1017), .in2(_42));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op312 (.out1(R313), .clock(clock), .in1(R312));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op439 (.out1(R440), .clock(clock), .in1(R439));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op565 (.out1(R566), .clock(clock), .in1(R565));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op683 (.out1(R684), .clock(clock), .in1(R683));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op800 (.out1(R801), .clock(clock), .in1(R800));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op909 (.out1(R910), .clock(clock), .in1(R909));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1017 (.out1(R1018), .clock(clock), .in1(idx_243));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op49 (.out1(_43), .in1(R1018));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op50 (.out1(_44), .in1(_43), .in2(2 'd 2));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op313 (.out1(R314), .clock(clock), .in1(R313));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op440 (.out1(R441), .clock(clock), .in1(R440));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op566 (.out1(R567), .clock(clock), .in1(R566));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op684 (.out1(R685), .clock(clock), .in1(R684));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op801 (.out1(R802), .clock(clock), .in1(R801));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op910 (.out1(R911), .clock(clock), .in1(R910));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1018 (.out1(R1019), .clock(clock), .in1(R1018));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op1118 (.out1(R1119), .clock(clock), .in1(_44));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op51 (.out1(_45), .in1(C40_244_D), .in2(R1119));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op314 (.out1(R315), .clock(clock), .in1(R314));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op441 (.out1(R442), .clock(clock), .in1(R441));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op567 (.out1(R568), .clock(clock), .in1(R567));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op685 (.out1(R686), .clock(clock), .in1(R685));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op802 (.out1(R803), .clock(clock), .in1(R802));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op911 (.out1(R912), .clock(clock), .in1(R911));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1019 (.out1(R1020), .clock(clock), .in1(R1019));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op1119 (.out1(R1120), .clock(clock), .in1(_45));
  SRAM op52 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_46),.ADR(R1120));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op315 (.out1(R316), .clock(clock), .in1(R315));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op442 (.out1(R443), .clock(clock), .in1(R442));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op568 (.out1(R569), .clock(clock), .in1(R568));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op686 (.out1(R687), .clock(clock), .in1(R686));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op803 (.out1(R804), .clock(clock), .in1(R803));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op912 (.out1(R913), .clock(clock), .in1(R912));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1020 (.out1(R1021), .clock(clock), .in1(R1020));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1120 (.out1(R1121), .clock(clock), .in1(_46));
  NE_EXPR #(.BITSIZE_in1(32), .BITSIZE_in2(1),.BITSIZE_out1(1)) op53 (.out1(ifout53), .in1(R1121), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op54 (.out1(_47), .in1(R1021));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op55 (.out1(_48), .in1(_47), .in2(2 'd 2));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op316 (.out1(R317), .clock(clock), .in1(R316));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op443 (.out1(R444), .clock(clock), .in1(R443));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op569 (.out1(R570), .clock(clock), .in1(R569));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op687 (.out1(R688), .clock(clock), .in1(R687));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op804 (.out1(R805), .clock(clock), .in1(R804));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op913 (.out1(R914), .clock(clock), .in1(R913));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1021 (.out1(R1022), .clock(clock), .in1(R1021));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1121 (.out1(R1122), .clock(clock), .in1(ifout53));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op1220 (.out1(R1221), .clock(clock), .in1(_48));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op56 (.out1(_49), .in1(C40_244_D), .in2(R1221));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op317 (.out1(R318), .clock(clock), .in1(R317));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op444 (.out1(R445), .clock(clock), .in1(R444));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op570 (.out1(R571), .clock(clock), .in1(R570));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op688 (.out1(R689), .clock(clock), .in1(R688));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op805 (.out1(R806), .clock(clock), .in1(R805));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op914 (.out1(R915), .clock(clock), .in1(R914));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1022 (.out1(R1023), .clock(clock), .in1(R1022));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1122 (.out1(R1123), .clock(clock), .in1(R1122));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op1221 (.out1(R1222), .clock(clock), .in1(_49));
  SRAM op57 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_50),.ADR(R1222));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op318 (.out1(R319), .clock(clock), .in1(R318));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op445 (.out1(R446), .clock(clock), .in1(R445));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op571 (.out1(R572), .clock(clock), .in1(R571));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op689 (.out1(R690), .clock(clock), .in1(R689));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op806 (.out1(R807), .clock(clock), .in1(R806));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op915 (.out1(R916), .clock(clock), .in1(R915));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1023 (.out1(R1024), .clock(clock), .in1(R1023));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1123 (.out1(R1124), .clock(clock), .in1(R1123));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1222 (.out1(R1223), .clock(clock), .in1(_50));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op58 (.out1(_51), .in1(R1223), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op319 (.out1(R320), .clock(clock), .in1(R319));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op446 (.out1(R447), .clock(clock), .in1(R446));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op572 (.out1(R573), .clock(clock), .in1(R572));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op690 (.out1(R691), .clock(clock), .in1(R690));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op807 (.out1(R808), .clock(clock), .in1(R807));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op916 (.out1(R917), .clock(clock), .in1(R916));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1024 (.out1(R1025), .clock(clock), .in1(R1024));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1124 (.out1(R1125), .clock(clock), .in1(R1124));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1223 (.out1(R1224), .clock(clock), .in1(_51));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(4), .BITSIZE_out1(32), .PRECISION(32)) op59 (.out1(_52), .in1(R1224), .in2(4 'd 8));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op320 (.out1(R321), .clock(clock), .in1(R320));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op447 (.out1(R448), .clock(clock), .in1(R447));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op573 (.out1(R574), .clock(clock), .in1(R573));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op691 (.out1(R692), .clock(clock), .in1(R691));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op808 (.out1(R809), .clock(clock), .in1(R808));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op917 (.out1(R918), .clock(clock), .in1(R917));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1025 (.out1(R1026), .clock(clock), .in1(R1025));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1125 (.out1(R1126), .clock(clock), .in1(R1125));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1224 (.out1(R1225), .clock(clock), .in1(_52));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(5), .BITSIZE_out1(64), .PRECISION(64)) op60 (.out1(_53), .in1(ip1_229_D), .in2(5 'd 16));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op61 (.out1(_54), .in1(_53));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(8), .BITSIZE_out1(32)) op62 (.out1(_55), .in1(_54), .in2(8 'd 255));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op63 (.out1(idx_247), .in1(R1225), .in2(_55));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op321 (.out1(R322), .clock(clock), .in1(R321));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op448 (.out1(R449), .clock(clock), .in1(R448));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op574 (.out1(R575), .clock(clock), .in1(R574));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op692 (.out1(R693), .clock(clock), .in1(R692));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op809 (.out1(R810), .clock(clock), .in1(R809));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op918 (.out1(R919), .clock(clock), .in1(R918));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1026 (.out1(R1027), .clock(clock), .in1(R1026));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1126 (.out1(R1127), .clock(clock), .in1(R1126));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1225 (.out1(R1226), .clock(clock), .in1(idx_247));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op64 (.out1(_56), .in1(R1226));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op65 (.out1(_57), .in1(_56), .in2(2 'd 2));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op322 (.out1(R323), .clock(clock), .in1(R322));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op449 (.out1(R450), .clock(clock), .in1(R449));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op575 (.out1(R576), .clock(clock), .in1(R575));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op693 (.out1(R694), .clock(clock), .in1(R693));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op810 (.out1(R811), .clock(clock), .in1(R810));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op919 (.out1(R920), .clock(clock), .in1(R919));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1027 (.out1(R1028), .clock(clock), .in1(R1027));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1127 (.out1(R1128), .clock(clock), .in1(R1127));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1226 (.out1(R1227), .clock(clock), .in1(R1226));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op1317 (.out1(R1318), .clock(clock), .in1(_57));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op66 (.out1(_58), .in1(C48_248_D), .in2(R1318));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op323 (.out1(R324), .clock(clock), .in1(R323));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op450 (.out1(R451), .clock(clock), .in1(R450));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op576 (.out1(R577), .clock(clock), .in1(R576));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op694 (.out1(R695), .clock(clock), .in1(R694));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op811 (.out1(R812), .clock(clock), .in1(R811));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op920 (.out1(R921), .clock(clock), .in1(R920));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1028 (.out1(R1029), .clock(clock), .in1(R1028));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1128 (.out1(R1129), .clock(clock), .in1(R1128));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1227 (.out1(R1228), .clock(clock), .in1(R1227));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op1318 (.out1(R1319), .clock(clock), .in1(_58));
  SRAM op67 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_59),.ADR(R1319));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op324 (.out1(R325), .clock(clock), .in1(R324));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op451 (.out1(R452), .clock(clock), .in1(R451));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op577 (.out1(R578), .clock(clock), .in1(R577));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op695 (.out1(R696), .clock(clock), .in1(R695));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op812 (.out1(R813), .clock(clock), .in1(R812));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op921 (.out1(R922), .clock(clock), .in1(R921));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1029 (.out1(R1030), .clock(clock), .in1(R1029));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1129 (.out1(R1130), .clock(clock), .in1(R1129));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1228 (.out1(R1229), .clock(clock), .in1(R1228));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1319 (.out1(R1320), .clock(clock), .in1(_59));
  NE_EXPR #(.BITSIZE_in1(32), .BITSIZE_in2(1),.BITSIZE_out1(1)) op68 (.out1(ifout68), .in1(R1320), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op69 (.out1(_60), .in1(R1229));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op70 (.out1(_61), .in1(_60), .in2(2 'd 2));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op325 (.out1(R326), .clock(clock), .in1(R325));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op452 (.out1(R453), .clock(clock), .in1(R452));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op578 (.out1(R579), .clock(clock), .in1(R578));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op696 (.out1(R697), .clock(clock), .in1(R696));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op813 (.out1(R814), .clock(clock), .in1(R813));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op922 (.out1(R923), .clock(clock), .in1(R922));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1030 (.out1(R1031), .clock(clock), .in1(R1030));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1130 (.out1(R1131), .clock(clock), .in1(R1130));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1229 (.out1(R1230), .clock(clock), .in1(R1229));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1320 (.out1(R1321), .clock(clock), .in1(ifout68));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op1410 (.out1(R1411), .clock(clock), .in1(_61));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op71 (.out1(_62), .in1(C48_248_D), .in2(R1411));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op326 (.out1(R327), .clock(clock), .in1(R326));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op453 (.out1(R454), .clock(clock), .in1(R453));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op579 (.out1(R580), .clock(clock), .in1(R579));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op697 (.out1(R698), .clock(clock), .in1(R697));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op814 (.out1(R815), .clock(clock), .in1(R814));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op923 (.out1(R924), .clock(clock), .in1(R923));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1031 (.out1(R1032), .clock(clock), .in1(R1031));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1131 (.out1(R1132), .clock(clock), .in1(R1131));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1230 (.out1(R1231), .clock(clock), .in1(R1230));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1321 (.out1(R1322), .clock(clock), .in1(R1321));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op1411 (.out1(R1412), .clock(clock), .in1(_62));
  SRAM op72 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_63),.ADR(R1412));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op327 (.out1(R328), .clock(clock), .in1(R327));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op454 (.out1(R455), .clock(clock), .in1(R454));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op580 (.out1(R581), .clock(clock), .in1(R580));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op698 (.out1(R699), .clock(clock), .in1(R698));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op815 (.out1(R816), .clock(clock), .in1(R815));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op924 (.out1(R925), .clock(clock), .in1(R924));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1032 (.out1(R1033), .clock(clock), .in1(R1032));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1132 (.out1(R1133), .clock(clock), .in1(R1132));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1231 (.out1(R1232), .clock(clock), .in1(R1231));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1322 (.out1(R1323), .clock(clock), .in1(R1322));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1412 (.out1(R1413), .clock(clock), .in1(_63));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op73 (.out1(_64), .in1(R1413), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op328 (.out1(R329), .clock(clock), .in1(R328));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op455 (.out1(R456), .clock(clock), .in1(R455));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op581 (.out1(R582), .clock(clock), .in1(R581));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op699 (.out1(R700), .clock(clock), .in1(R699));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op816 (.out1(R817), .clock(clock), .in1(R816));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op925 (.out1(R926), .clock(clock), .in1(R925));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1033 (.out1(R1034), .clock(clock), .in1(R1033));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1133 (.out1(R1134), .clock(clock), .in1(R1133));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1232 (.out1(R1233), .clock(clock), .in1(R1232));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1323 (.out1(R1324), .clock(clock), .in1(R1323));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1413 (.out1(R1414), .clock(clock), .in1(_64));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(4), .BITSIZE_out1(32), .PRECISION(32)) op74 (.out1(_65), .in1(R1414), .in2(4 'd 8));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op329 (.out1(R330), .clock(clock), .in1(R329));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op456 (.out1(R457), .clock(clock), .in1(R456));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op582 (.out1(R583), .clock(clock), .in1(R582));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op700 (.out1(R701), .clock(clock), .in1(R700));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op817 (.out1(R818), .clock(clock), .in1(R817));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op926 (.out1(R927), .clock(clock), .in1(R926));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1034 (.out1(R1035), .clock(clock), .in1(R1034));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1134 (.out1(R1135), .clock(clock), .in1(R1134));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1233 (.out1(R1234), .clock(clock), .in1(R1233));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1324 (.out1(R1325), .clock(clock), .in1(R1324));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1414 (.out1(R1415), .clock(clock), .in1(_65));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(4), .BITSIZE_out1(64), .PRECISION(64)) op75 (.out1(_66), .in1(ip1_229_D), .in2(4 'd 8));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op76 (.out1(_67), .in1(_66));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(8), .BITSIZE_out1(32)) op77 (.out1(_68), .in1(_67), .in2(8 'd 255));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op78 (.out1(idx_251), .in1(R1415), .in2(_68));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op330 (.out1(R331), .clock(clock), .in1(R330));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op457 (.out1(R458), .clock(clock), .in1(R457));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op583 (.out1(R584), .clock(clock), .in1(R583));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op701 (.out1(R702), .clock(clock), .in1(R701));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op818 (.out1(R819), .clock(clock), .in1(R818));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op927 (.out1(R928), .clock(clock), .in1(R927));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1035 (.out1(R1036), .clock(clock), .in1(R1035));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1135 (.out1(R1136), .clock(clock), .in1(R1135));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1234 (.out1(R1235), .clock(clock), .in1(R1234));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1325 (.out1(R1326), .clock(clock), .in1(R1325));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1415 (.out1(R1416), .clock(clock), .in1(idx_251));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op79 (.out1(_69), .in1(R1416));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op80 (.out1(_70), .in1(_69), .in2(2 'd 2));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op331 (.out1(R332), .clock(clock), .in1(R331));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op458 (.out1(R459), .clock(clock), .in1(R458));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op584 (.out1(R585), .clock(clock), .in1(R584));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op702 (.out1(R703), .clock(clock), .in1(R702));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op819 (.out1(R820), .clock(clock), .in1(R819));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op928 (.out1(R929), .clock(clock), .in1(R928));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1036 (.out1(R1037), .clock(clock), .in1(R1036));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1136 (.out1(R1137), .clock(clock), .in1(R1136));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1235 (.out1(R1236), .clock(clock), .in1(R1235));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1326 (.out1(R1327), .clock(clock), .in1(R1326));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1416 (.out1(R1417), .clock(clock), .in1(R1416));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op1498 (.out1(R1499), .clock(clock), .in1(_70));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op81 (.out1(_71), .in1(C56_252_D), .in2(R1499));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op332 (.out1(R333), .clock(clock), .in1(R332));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op459 (.out1(R460), .clock(clock), .in1(R459));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op585 (.out1(R586), .clock(clock), .in1(R585));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op703 (.out1(R704), .clock(clock), .in1(R703));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op820 (.out1(R821), .clock(clock), .in1(R820));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op929 (.out1(R930), .clock(clock), .in1(R929));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1037 (.out1(R1038), .clock(clock), .in1(R1037));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1137 (.out1(R1138), .clock(clock), .in1(R1137));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1236 (.out1(R1237), .clock(clock), .in1(R1236));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1327 (.out1(R1328), .clock(clock), .in1(R1327));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1417 (.out1(R1418), .clock(clock), .in1(R1417));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op1499 (.out1(R1500), .clock(clock), .in1(_71));
  SRAM op82 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_72),.ADR(R1500));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op333 (.out1(R334), .clock(clock), .in1(R333));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op460 (.out1(R461), .clock(clock), .in1(R460));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op586 (.out1(R587), .clock(clock), .in1(R586));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op704 (.out1(R705), .clock(clock), .in1(R704));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op821 (.out1(R822), .clock(clock), .in1(R821));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op930 (.out1(R931), .clock(clock), .in1(R930));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1038 (.out1(R1039), .clock(clock), .in1(R1038));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1138 (.out1(R1139), .clock(clock), .in1(R1138));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1237 (.out1(R1238), .clock(clock), .in1(R1237));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1328 (.out1(R1329), .clock(clock), .in1(R1328));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1418 (.out1(R1419), .clock(clock), .in1(R1418));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1500 (.out1(R1501), .clock(clock), .in1(_72));
  NE_EXPR #(.BITSIZE_in1(32), .BITSIZE_in2(1),.BITSIZE_out1(1)) op83 (.out1(ifout83), .in1(R1501), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op84 (.out1(_73), .in1(R1419));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op85 (.out1(_74), .in1(_73), .in2(2 'd 2));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op334 (.out1(R335), .clock(clock), .in1(R334));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op461 (.out1(R462), .clock(clock), .in1(R461));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op587 (.out1(R588), .clock(clock), .in1(R587));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op705 (.out1(R706), .clock(clock), .in1(R705));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op822 (.out1(R823), .clock(clock), .in1(R822));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op931 (.out1(R932), .clock(clock), .in1(R931));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1039 (.out1(R1040), .clock(clock), .in1(R1039));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1139 (.out1(R1140), .clock(clock), .in1(R1139));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1238 (.out1(R1239), .clock(clock), .in1(R1238));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1329 (.out1(R1330), .clock(clock), .in1(R1329));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1419 (.out1(R1420), .clock(clock), .in1(R1419));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1501 (.out1(R1502), .clock(clock), .in1(ifout83));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op1582 (.out1(R1583), .clock(clock), .in1(_74));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op86 (.out1(_75), .in1(C56_252_D), .in2(R1583));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op335 (.out1(R336), .clock(clock), .in1(R335));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op462 (.out1(R463), .clock(clock), .in1(R462));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op588 (.out1(R589), .clock(clock), .in1(R588));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op706 (.out1(R707), .clock(clock), .in1(R706));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op823 (.out1(R824), .clock(clock), .in1(R823));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op932 (.out1(R933), .clock(clock), .in1(R932));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1040 (.out1(R1041), .clock(clock), .in1(R1040));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1140 (.out1(R1141), .clock(clock), .in1(R1140));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1239 (.out1(R1240), .clock(clock), .in1(R1239));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1330 (.out1(R1331), .clock(clock), .in1(R1330));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1420 (.out1(R1421), .clock(clock), .in1(R1420));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1502 (.out1(R1503), .clock(clock), .in1(R1502));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op1583 (.out1(R1584), .clock(clock), .in1(_75));
  SRAM op87 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_76),.ADR(R1584));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op336 (.out1(R337), .clock(clock), .in1(R336));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op463 (.out1(R464), .clock(clock), .in1(R463));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op589 (.out1(R590), .clock(clock), .in1(R589));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op707 (.out1(R708), .clock(clock), .in1(R707));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op824 (.out1(R825), .clock(clock), .in1(R824));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op933 (.out1(R934), .clock(clock), .in1(R933));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1041 (.out1(R1042), .clock(clock), .in1(R1041));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1141 (.out1(R1142), .clock(clock), .in1(R1141));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1240 (.out1(R1241), .clock(clock), .in1(R1240));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1331 (.out1(R1332), .clock(clock), .in1(R1331));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1421 (.out1(R1422), .clock(clock), .in1(R1421));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1503 (.out1(R1504), .clock(clock), .in1(R1503));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1584 (.out1(R1585), .clock(clock), .in1(_76));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op88 (.out1(_77), .in1(R1585), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op337 (.out1(R338), .clock(clock), .in1(R337));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op464 (.out1(R465), .clock(clock), .in1(R464));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op590 (.out1(R591), .clock(clock), .in1(R590));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op708 (.out1(R709), .clock(clock), .in1(R708));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op825 (.out1(R826), .clock(clock), .in1(R825));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op934 (.out1(R935), .clock(clock), .in1(R934));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1042 (.out1(R1043), .clock(clock), .in1(R1042));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1142 (.out1(R1143), .clock(clock), .in1(R1142));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1241 (.out1(R1242), .clock(clock), .in1(R1241));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1332 (.out1(R1333), .clock(clock), .in1(R1332));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1422 (.out1(R1423), .clock(clock), .in1(R1422));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1504 (.out1(R1505), .clock(clock), .in1(R1504));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1585 (.out1(R1586), .clock(clock), .in1(_77));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(4), .BITSIZE_out1(32), .PRECISION(32)) op89 (.out1(_78), .in1(R1586), .in2(4 'd 8));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op338 (.out1(R339), .clock(clock), .in1(R338));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op465 (.out1(R466), .clock(clock), .in1(R465));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op591 (.out1(R592), .clock(clock), .in1(R591));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op709 (.out1(R710), .clock(clock), .in1(R709));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op826 (.out1(R827), .clock(clock), .in1(R826));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op935 (.out1(R936), .clock(clock), .in1(R935));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1043 (.out1(R1044), .clock(clock), .in1(R1043));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1143 (.out1(R1144), .clock(clock), .in1(R1143));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1242 (.out1(R1243), .clock(clock), .in1(R1242));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1333 (.out1(R1334), .clock(clock), .in1(R1333));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1423 (.out1(R1424), .clock(clock), .in1(R1423));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1505 (.out1(R1506), .clock(clock), .in1(R1505));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1586 (.out1(R1587), .clock(clock), .in1(_78));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op90 (.out1(_79), .in1(ip1_229_D));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(8), .BITSIZE_out1(32)) op91 (.out1(_80), .in1(_79), .in2(8 'd 255));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op92 (.out1(idx_255), .in1(R1587), .in2(_80));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op339 (.out1(R340), .clock(clock), .in1(R339));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op466 (.out1(R467), .clock(clock), .in1(R466));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op592 (.out1(R593), .clock(clock), .in1(R592));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op710 (.out1(R711), .clock(clock), .in1(R710));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op827 (.out1(R828), .clock(clock), .in1(R827));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op936 (.out1(R937), .clock(clock), .in1(R936));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1044 (.out1(R1045), .clock(clock), .in1(R1044));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1144 (.out1(R1145), .clock(clock), .in1(R1144));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1243 (.out1(R1244), .clock(clock), .in1(R1243));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1334 (.out1(R1335), .clock(clock), .in1(R1334));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1424 (.out1(R1425), .clock(clock), .in1(R1424));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1506 (.out1(R1507), .clock(clock), .in1(R1506));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1587 (.out1(R1588), .clock(clock), .in1(idx_255));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op93 (.out1(_81), .in1(R1588));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op94 (.out1(_82), .in1(_81), .in2(2 'd 2));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op340 (.out1(R341), .clock(clock), .in1(R340));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op467 (.out1(R468), .clock(clock), .in1(R467));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op593 (.out1(R594), .clock(clock), .in1(R593));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op711 (.out1(R712), .clock(clock), .in1(R711));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op828 (.out1(R829), .clock(clock), .in1(R828));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op937 (.out1(R938), .clock(clock), .in1(R937));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1045 (.out1(R1046), .clock(clock), .in1(R1045));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1145 (.out1(R1146), .clock(clock), .in1(R1145));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1244 (.out1(R1245), .clock(clock), .in1(R1244));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1335 (.out1(R1336), .clock(clock), .in1(R1335));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1425 (.out1(R1426), .clock(clock), .in1(R1425));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1507 (.out1(R1508), .clock(clock), .in1(R1507));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1588 (.out1(R1589), .clock(clock), .in1(R1588));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op1660 (.out1(R1661), .clock(clock), .in1(_82));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op95 (.out1(_83), .in1(C64_256_D), .in2(R1661));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op341 (.out1(R342), .clock(clock), .in1(R341));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op468 (.out1(R469), .clock(clock), .in1(R468));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op594 (.out1(R595), .clock(clock), .in1(R594));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op712 (.out1(R713), .clock(clock), .in1(R712));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op829 (.out1(R830), .clock(clock), .in1(R829));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op938 (.out1(R939), .clock(clock), .in1(R938));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1046 (.out1(R1047), .clock(clock), .in1(R1046));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1146 (.out1(R1147), .clock(clock), .in1(R1146));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1245 (.out1(R1246), .clock(clock), .in1(R1245));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1336 (.out1(R1337), .clock(clock), .in1(R1336));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1426 (.out1(R1427), .clock(clock), .in1(R1426));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1508 (.out1(R1509), .clock(clock), .in1(R1508));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1589 (.out1(R1590), .clock(clock), .in1(R1589));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op1661 (.out1(R1662), .clock(clock), .in1(_83));
  SRAM op96 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_84),.ADR(R1662));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op342 (.out1(R343), .clock(clock), .in1(R342));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op469 (.out1(R470), .clock(clock), .in1(R469));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op595 (.out1(R596), .clock(clock), .in1(R595));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op713 (.out1(R714), .clock(clock), .in1(R713));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op830 (.out1(R831), .clock(clock), .in1(R830));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op939 (.out1(R940), .clock(clock), .in1(R939));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1047 (.out1(R1048), .clock(clock), .in1(R1047));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1147 (.out1(R1148), .clock(clock), .in1(R1147));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1246 (.out1(R1247), .clock(clock), .in1(R1246));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1337 (.out1(R1338), .clock(clock), .in1(R1337));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1427 (.out1(R1428), .clock(clock), .in1(R1427));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1509 (.out1(R1510), .clock(clock), .in1(R1509));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1590 (.out1(R1591), .clock(clock), .in1(R1590));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1662 (.out1(R1663), .clock(clock), .in1(_84));
  NE_EXPR #(.BITSIZE_in1(32), .BITSIZE_in2(1),.BITSIZE_out1(1)) op97 (.out1(ifout97), .in1(R1663), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op98 (.out1(_85), .in1(R1591));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op99 (.out1(_86), .in1(_85), .in2(2 'd 2));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op343 (.out1(R344), .clock(clock), .in1(R343));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op470 (.out1(R471), .clock(clock), .in1(R470));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op596 (.out1(R597), .clock(clock), .in1(R596));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op714 (.out1(R715), .clock(clock), .in1(R714));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op831 (.out1(R832), .clock(clock), .in1(R831));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op940 (.out1(R941), .clock(clock), .in1(R940));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1048 (.out1(R1049), .clock(clock), .in1(R1048));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1148 (.out1(R1149), .clock(clock), .in1(R1148));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1247 (.out1(R1248), .clock(clock), .in1(R1247));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1338 (.out1(R1339), .clock(clock), .in1(R1338));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1428 (.out1(R1429), .clock(clock), .in1(R1428));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1510 (.out1(R1511), .clock(clock), .in1(R1510));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1591 (.out1(R1592), .clock(clock), .in1(R1591));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1663 (.out1(R1664), .clock(clock), .in1(ifout97));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op1735 (.out1(R1736), .clock(clock), .in1(_86));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op100 (.out1(_87), .in1(C64_256_D), .in2(R1736));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op344 (.out1(R345), .clock(clock), .in1(R344));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op471 (.out1(R472), .clock(clock), .in1(R471));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op597 (.out1(R598), .clock(clock), .in1(R597));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op715 (.out1(R716), .clock(clock), .in1(R715));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op832 (.out1(R833), .clock(clock), .in1(R832));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op941 (.out1(R942), .clock(clock), .in1(R941));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1049 (.out1(R1050), .clock(clock), .in1(R1049));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1149 (.out1(R1150), .clock(clock), .in1(R1149));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1248 (.out1(R1249), .clock(clock), .in1(R1248));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1339 (.out1(R1340), .clock(clock), .in1(R1339));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1429 (.out1(R1430), .clock(clock), .in1(R1429));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1511 (.out1(R1512), .clock(clock), .in1(R1511));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1592 (.out1(R1593), .clock(clock), .in1(R1592));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1664 (.out1(R1665), .clock(clock), .in1(R1664));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op1736 (.out1(R1737), .clock(clock), .in1(_87));
  SRAM op101 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_88),.ADR(R1737));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op345 (.out1(R346), .clock(clock), .in1(R345));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op472 (.out1(R473), .clock(clock), .in1(R472));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op598 (.out1(R599), .clock(clock), .in1(R598));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op716 (.out1(R717), .clock(clock), .in1(R716));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op833 (.out1(R834), .clock(clock), .in1(R833));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op942 (.out1(R943), .clock(clock), .in1(R942));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1050 (.out1(R1051), .clock(clock), .in1(R1050));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1150 (.out1(R1151), .clock(clock), .in1(R1150));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1249 (.out1(R1250), .clock(clock), .in1(R1249));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1340 (.out1(R1341), .clock(clock), .in1(R1340));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1430 (.out1(R1431), .clock(clock), .in1(R1430));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1512 (.out1(R1513), .clock(clock), .in1(R1512));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1593 (.out1(R1594), .clock(clock), .in1(R1593));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1665 (.out1(R1666), .clock(clock), .in1(R1665));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1737 (.out1(R1738), .clock(clock), .in1(_88));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op102 (.out1(_89), .in1(R1738), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op346 (.out1(R347), .clock(clock), .in1(R346));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op473 (.out1(R474), .clock(clock), .in1(R473));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op599 (.out1(R600), .clock(clock), .in1(R599));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op717 (.out1(R718), .clock(clock), .in1(R717));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op834 (.out1(R835), .clock(clock), .in1(R834));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op943 (.out1(R944), .clock(clock), .in1(R943));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1051 (.out1(R1052), .clock(clock), .in1(R1051));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1151 (.out1(R1152), .clock(clock), .in1(R1151));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1250 (.out1(R1251), .clock(clock), .in1(R1250));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1341 (.out1(R1342), .clock(clock), .in1(R1341));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1431 (.out1(R1432), .clock(clock), .in1(R1431));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1513 (.out1(R1514), .clock(clock), .in1(R1513));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1594 (.out1(R1595), .clock(clock), .in1(R1594));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1666 (.out1(R1667), .clock(clock), .in1(R1666));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1738 (.out1(R1739), .clock(clock), .in1(_89));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(4), .BITSIZE_out1(32), .PRECISION(32)) op103 (.out1(_90), .in1(R1739), .in2(4 'd 8));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op347 (.out1(R348), .clock(clock), .in1(R347));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op474 (.out1(R475), .clock(clock), .in1(R474));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op600 (.out1(R601), .clock(clock), .in1(R600));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op718 (.out1(R719), .clock(clock), .in1(R718));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op835 (.out1(R836), .clock(clock), .in1(R835));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op944 (.out1(R945), .clock(clock), .in1(R944));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1052 (.out1(R1053), .clock(clock), .in1(R1052));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1152 (.out1(R1153), .clock(clock), .in1(R1152));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1251 (.out1(R1252), .clock(clock), .in1(R1251));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1342 (.out1(R1343), .clock(clock), .in1(R1342));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1432 (.out1(R1433), .clock(clock), .in1(R1432));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1514 (.out1(R1515), .clock(clock), .in1(R1514));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1595 (.out1(R1596), .clock(clock), .in1(R1595));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1667 (.out1(R1668), .clock(clock), .in1(R1667));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1739 (.out1(R1740), .clock(clock), .in1(_90));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op104 (.out1(_91), .in1(ip2_259_D), .in2(6 'd 56));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op105 (.out1(_92), .in1(_91));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op106 (.out1(idx_260), .in1(R1740), .in2(_92));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op348 (.out1(R349), .clock(clock), .in1(R348));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op475 (.out1(R476), .clock(clock), .in1(R475));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op601 (.out1(R602), .clock(clock), .in1(R601));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op719 (.out1(R720), .clock(clock), .in1(R719));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op836 (.out1(R837), .clock(clock), .in1(R836));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op945 (.out1(R946), .clock(clock), .in1(R945));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1053 (.out1(R1054), .clock(clock), .in1(R1053));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1153 (.out1(R1154), .clock(clock), .in1(R1153));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1252 (.out1(R1253), .clock(clock), .in1(R1252));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1343 (.out1(R1344), .clock(clock), .in1(R1343));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1433 (.out1(R1434), .clock(clock), .in1(R1433));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1515 (.out1(R1516), .clock(clock), .in1(R1515));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1596 (.out1(R1597), .clock(clock), .in1(R1596));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1668 (.out1(R1669), .clock(clock), .in1(R1668));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1740 (.out1(R1741), .clock(clock), .in1(idx_260));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op107 (.out1(_93), .in1(R1741));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op108 (.out1(_94), .in1(_93), .in2(2 'd 2));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op349 (.out1(R350), .clock(clock), .in1(R349));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op476 (.out1(R477), .clock(clock), .in1(R476));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op602 (.out1(R603), .clock(clock), .in1(R602));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op720 (.out1(R721), .clock(clock), .in1(R720));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op837 (.out1(R838), .clock(clock), .in1(R837));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op946 (.out1(R947), .clock(clock), .in1(R946));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1054 (.out1(R1055), .clock(clock), .in1(R1054));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1154 (.out1(R1155), .clock(clock), .in1(R1154));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1253 (.out1(R1254), .clock(clock), .in1(R1253));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1344 (.out1(R1345), .clock(clock), .in1(R1344));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1434 (.out1(R1435), .clock(clock), .in1(R1434));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1516 (.out1(R1517), .clock(clock), .in1(R1516));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1597 (.out1(R1598), .clock(clock), .in1(R1597));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1669 (.out1(R1670), .clock(clock), .in1(R1669));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1741 (.out1(R1742), .clock(clock), .in1(R1741));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op1804 (.out1(R1805), .clock(clock), .in1(_94));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op109 (.out1(_95), .in1(C72_261_D), .in2(R1805));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op350 (.out1(R351), .clock(clock), .in1(R350));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op477 (.out1(R478), .clock(clock), .in1(R477));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op603 (.out1(R604), .clock(clock), .in1(R603));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op721 (.out1(R722), .clock(clock), .in1(R721));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op838 (.out1(R839), .clock(clock), .in1(R838));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op947 (.out1(R948), .clock(clock), .in1(R947));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1055 (.out1(R1056), .clock(clock), .in1(R1055));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1155 (.out1(R1156), .clock(clock), .in1(R1155));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1254 (.out1(R1255), .clock(clock), .in1(R1254));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1345 (.out1(R1346), .clock(clock), .in1(R1345));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1435 (.out1(R1436), .clock(clock), .in1(R1435));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1517 (.out1(R1518), .clock(clock), .in1(R1517));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1598 (.out1(R1599), .clock(clock), .in1(R1598));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1670 (.out1(R1671), .clock(clock), .in1(R1670));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1742 (.out1(R1743), .clock(clock), .in1(R1742));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op1805 (.out1(R1806), .clock(clock), .in1(_95));
  SRAM op110 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_96),.ADR(R1806));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op351 (.out1(R352), .clock(clock), .in1(R351));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op478 (.out1(R479), .clock(clock), .in1(R478));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op604 (.out1(R605), .clock(clock), .in1(R604));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op722 (.out1(R723), .clock(clock), .in1(R722));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op839 (.out1(R840), .clock(clock), .in1(R839));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op948 (.out1(R949), .clock(clock), .in1(R948));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1056 (.out1(R1057), .clock(clock), .in1(R1056));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1156 (.out1(R1157), .clock(clock), .in1(R1156));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1255 (.out1(R1256), .clock(clock), .in1(R1255));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1346 (.out1(R1347), .clock(clock), .in1(R1346));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1436 (.out1(R1437), .clock(clock), .in1(R1436));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1518 (.out1(R1519), .clock(clock), .in1(R1518));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1599 (.out1(R1600), .clock(clock), .in1(R1599));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1671 (.out1(R1672), .clock(clock), .in1(R1671));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1743 (.out1(R1744), .clock(clock), .in1(R1743));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1806 (.out1(R1807), .clock(clock), .in1(_96));
  NE_EXPR #(.BITSIZE_in1(32), .BITSIZE_in2(1),.BITSIZE_out1(1)) op111 (.out1(ifout111), .in1(R1807), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op112 (.out1(_97), .in1(R1744));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op113 (.out1(_98), .in1(_97), .in2(2 'd 2));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op352 (.out1(R353), .clock(clock), .in1(R352));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op479 (.out1(R480), .clock(clock), .in1(R479));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op605 (.out1(R606), .clock(clock), .in1(R605));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op723 (.out1(R724), .clock(clock), .in1(R723));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op840 (.out1(R841), .clock(clock), .in1(R840));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op949 (.out1(R950), .clock(clock), .in1(R949));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1057 (.out1(R1058), .clock(clock), .in1(R1057));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1157 (.out1(R1158), .clock(clock), .in1(R1157));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1256 (.out1(R1257), .clock(clock), .in1(R1256));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1347 (.out1(R1348), .clock(clock), .in1(R1347));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1437 (.out1(R1438), .clock(clock), .in1(R1437));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1519 (.out1(R1520), .clock(clock), .in1(R1519));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1600 (.out1(R1601), .clock(clock), .in1(R1600));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1672 (.out1(R1673), .clock(clock), .in1(R1672));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1744 (.out1(R1745), .clock(clock), .in1(R1744));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1807 (.out1(R1808), .clock(clock), .in1(ifout111));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op1870 (.out1(R1871), .clock(clock), .in1(_98));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op114 (.out1(_99), .in1(C72_261_D), .in2(R1871));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op353 (.out1(R354), .clock(clock), .in1(R353));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op480 (.out1(R481), .clock(clock), .in1(R480));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op606 (.out1(R607), .clock(clock), .in1(R606));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op724 (.out1(R725), .clock(clock), .in1(R724));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op841 (.out1(R842), .clock(clock), .in1(R841));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op950 (.out1(R951), .clock(clock), .in1(R950));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1058 (.out1(R1059), .clock(clock), .in1(R1058));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1158 (.out1(R1159), .clock(clock), .in1(R1158));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1257 (.out1(R1258), .clock(clock), .in1(R1257));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1348 (.out1(R1349), .clock(clock), .in1(R1348));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1438 (.out1(R1439), .clock(clock), .in1(R1438));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1520 (.out1(R1521), .clock(clock), .in1(R1520));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1601 (.out1(R1602), .clock(clock), .in1(R1601));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1673 (.out1(R1674), .clock(clock), .in1(R1673));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1745 (.out1(R1746), .clock(clock), .in1(R1745));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1808 (.out1(R1809), .clock(clock), .in1(R1808));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op1871 (.out1(R1872), .clock(clock), .in1(_99));
  SRAM op115 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_100),.ADR(R1872));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op354 (.out1(R355), .clock(clock), .in1(R354));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op481 (.out1(R482), .clock(clock), .in1(R481));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op607 (.out1(R608), .clock(clock), .in1(R607));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op725 (.out1(R726), .clock(clock), .in1(R725));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op842 (.out1(R843), .clock(clock), .in1(R842));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op951 (.out1(R952), .clock(clock), .in1(R951));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1059 (.out1(R1060), .clock(clock), .in1(R1059));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1159 (.out1(R1160), .clock(clock), .in1(R1159));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1258 (.out1(R1259), .clock(clock), .in1(R1258));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1349 (.out1(R1350), .clock(clock), .in1(R1349));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1439 (.out1(R1440), .clock(clock), .in1(R1439));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1521 (.out1(R1522), .clock(clock), .in1(R1521));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1602 (.out1(R1603), .clock(clock), .in1(R1602));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1674 (.out1(R1675), .clock(clock), .in1(R1674));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1746 (.out1(R1747), .clock(clock), .in1(R1746));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1809 (.out1(R1810), .clock(clock), .in1(R1809));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1872 (.out1(R1873), .clock(clock), .in1(_100));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op116 (.out1(_101), .in1(R1873), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op355 (.out1(R356), .clock(clock), .in1(R355));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op482 (.out1(R483), .clock(clock), .in1(R482));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op608 (.out1(R609), .clock(clock), .in1(R608));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op726 (.out1(R727), .clock(clock), .in1(R726));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op843 (.out1(R844), .clock(clock), .in1(R843));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op952 (.out1(R953), .clock(clock), .in1(R952));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1060 (.out1(R1061), .clock(clock), .in1(R1060));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1160 (.out1(R1161), .clock(clock), .in1(R1160));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1259 (.out1(R1260), .clock(clock), .in1(R1259));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1350 (.out1(R1351), .clock(clock), .in1(R1350));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1440 (.out1(R1441), .clock(clock), .in1(R1440));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1522 (.out1(R1523), .clock(clock), .in1(R1522));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1603 (.out1(R1604), .clock(clock), .in1(R1603));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1675 (.out1(R1676), .clock(clock), .in1(R1675));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1747 (.out1(R1748), .clock(clock), .in1(R1747));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1810 (.out1(R1811), .clock(clock), .in1(R1810));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1873 (.out1(R1874), .clock(clock), .in1(_101));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(4), .BITSIZE_out1(32), .PRECISION(32)) op117 (.out1(_102), .in1(R1874), .in2(4 'd 8));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op356 (.out1(R357), .clock(clock), .in1(R356));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op483 (.out1(R484), .clock(clock), .in1(R483));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op609 (.out1(R610), .clock(clock), .in1(R609));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op727 (.out1(R728), .clock(clock), .in1(R727));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op844 (.out1(R845), .clock(clock), .in1(R844));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op953 (.out1(R954), .clock(clock), .in1(R953));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1061 (.out1(R1062), .clock(clock), .in1(R1061));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1161 (.out1(R1162), .clock(clock), .in1(R1161));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1260 (.out1(R1261), .clock(clock), .in1(R1260));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1351 (.out1(R1352), .clock(clock), .in1(R1351));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1441 (.out1(R1442), .clock(clock), .in1(R1441));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1523 (.out1(R1524), .clock(clock), .in1(R1523));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1604 (.out1(R1605), .clock(clock), .in1(R1604));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1676 (.out1(R1677), .clock(clock), .in1(R1676));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1748 (.out1(R1749), .clock(clock), .in1(R1748));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1811 (.out1(R1812), .clock(clock), .in1(R1811));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1874 (.out1(R1875), .clock(clock), .in1(_102));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op118 (.out1(_103), .in1(ip2_259_D), .in2(6 'd 48));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op119 (.out1(_104), .in1(_103));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(8), .BITSIZE_out1(32)) op120 (.out1(_105), .in1(_104), .in2(8 'd 255));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op121 (.out1(idx_264), .in1(R1875), .in2(_105));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op357 (.out1(R358), .clock(clock), .in1(R357));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op484 (.out1(R485), .clock(clock), .in1(R484));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op610 (.out1(R611), .clock(clock), .in1(R610));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op728 (.out1(R729), .clock(clock), .in1(R728));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op845 (.out1(R846), .clock(clock), .in1(R845));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op954 (.out1(R955), .clock(clock), .in1(R954));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1062 (.out1(R1063), .clock(clock), .in1(R1062));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1162 (.out1(R1163), .clock(clock), .in1(R1162));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1261 (.out1(R1262), .clock(clock), .in1(R1261));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1352 (.out1(R1353), .clock(clock), .in1(R1352));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1442 (.out1(R1443), .clock(clock), .in1(R1442));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1524 (.out1(R1525), .clock(clock), .in1(R1524));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1605 (.out1(R1606), .clock(clock), .in1(R1605));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1677 (.out1(R1678), .clock(clock), .in1(R1677));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1749 (.out1(R1750), .clock(clock), .in1(R1749));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1812 (.out1(R1813), .clock(clock), .in1(R1812));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1875 (.out1(R1876), .clock(clock), .in1(idx_264));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op122 (.out1(_106), .in1(R1876));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op123 (.out1(_107), .in1(_106), .in2(2 'd 2));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op358 (.out1(R359), .clock(clock), .in1(R358));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op485 (.out1(R486), .clock(clock), .in1(R485));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op611 (.out1(R612), .clock(clock), .in1(R611));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op729 (.out1(R730), .clock(clock), .in1(R729));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op846 (.out1(R847), .clock(clock), .in1(R846));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op955 (.out1(R956), .clock(clock), .in1(R955));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1063 (.out1(R1064), .clock(clock), .in1(R1063));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1163 (.out1(R1164), .clock(clock), .in1(R1163));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1262 (.out1(R1263), .clock(clock), .in1(R1262));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1353 (.out1(R1354), .clock(clock), .in1(R1353));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1443 (.out1(R1444), .clock(clock), .in1(R1443));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1525 (.out1(R1526), .clock(clock), .in1(R1525));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1606 (.out1(R1607), .clock(clock), .in1(R1606));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1678 (.out1(R1679), .clock(clock), .in1(R1678));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1750 (.out1(R1751), .clock(clock), .in1(R1750));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1813 (.out1(R1814), .clock(clock), .in1(R1813));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1876 (.out1(R1877), .clock(clock), .in1(R1876));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op1930 (.out1(R1931), .clock(clock), .in1(_107));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op124 (.out1(_108), .in1(C80_265_D), .in2(R1931));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op359 (.out1(R360), .clock(clock), .in1(R359));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op486 (.out1(R487), .clock(clock), .in1(R486));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op612 (.out1(R613), .clock(clock), .in1(R612));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op730 (.out1(R731), .clock(clock), .in1(R730));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op847 (.out1(R848), .clock(clock), .in1(R847));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op956 (.out1(R957), .clock(clock), .in1(R956));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1064 (.out1(R1065), .clock(clock), .in1(R1064));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1164 (.out1(R1165), .clock(clock), .in1(R1164));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1263 (.out1(R1264), .clock(clock), .in1(R1263));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1354 (.out1(R1355), .clock(clock), .in1(R1354));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1444 (.out1(R1445), .clock(clock), .in1(R1444));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1526 (.out1(R1527), .clock(clock), .in1(R1526));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1607 (.out1(R1608), .clock(clock), .in1(R1607));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1679 (.out1(R1680), .clock(clock), .in1(R1679));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1751 (.out1(R1752), .clock(clock), .in1(R1751));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1814 (.out1(R1815), .clock(clock), .in1(R1814));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1877 (.out1(R1878), .clock(clock), .in1(R1877));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op1931 (.out1(R1932), .clock(clock), .in1(_108));
  SRAM op125 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_109),.ADR(R1932));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op360 (.out1(R361), .clock(clock), .in1(R360));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op487 (.out1(R488), .clock(clock), .in1(R487));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op613 (.out1(R614), .clock(clock), .in1(R613));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op731 (.out1(R732), .clock(clock), .in1(R731));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op848 (.out1(R849), .clock(clock), .in1(R848));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op957 (.out1(R958), .clock(clock), .in1(R957));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1065 (.out1(R1066), .clock(clock), .in1(R1065));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1165 (.out1(R1166), .clock(clock), .in1(R1165));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1264 (.out1(R1265), .clock(clock), .in1(R1264));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1355 (.out1(R1356), .clock(clock), .in1(R1355));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1445 (.out1(R1446), .clock(clock), .in1(R1445));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1527 (.out1(R1528), .clock(clock), .in1(R1527));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1608 (.out1(R1609), .clock(clock), .in1(R1608));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1680 (.out1(R1681), .clock(clock), .in1(R1680));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1752 (.out1(R1753), .clock(clock), .in1(R1752));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1815 (.out1(R1816), .clock(clock), .in1(R1815));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1878 (.out1(R1879), .clock(clock), .in1(R1878));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1932 (.out1(R1933), .clock(clock), .in1(_109));
  NE_EXPR #(.BITSIZE_in1(32), .BITSIZE_in2(1),.BITSIZE_out1(1)) op126 (.out1(ifout126), .in1(R1933), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op127 (.out1(_110), .in1(R1879));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op128 (.out1(_111), .in1(_110), .in2(2 'd 2));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op361 (.out1(R362), .clock(clock), .in1(R361));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op488 (.out1(R489), .clock(clock), .in1(R488));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op614 (.out1(R615), .clock(clock), .in1(R614));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op732 (.out1(R733), .clock(clock), .in1(R732));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op849 (.out1(R850), .clock(clock), .in1(R849));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op958 (.out1(R959), .clock(clock), .in1(R958));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1066 (.out1(R1067), .clock(clock), .in1(R1066));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1166 (.out1(R1167), .clock(clock), .in1(R1166));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1265 (.out1(R1266), .clock(clock), .in1(R1265));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1356 (.out1(R1357), .clock(clock), .in1(R1356));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1446 (.out1(R1447), .clock(clock), .in1(R1446));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1528 (.out1(R1529), .clock(clock), .in1(R1528));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1609 (.out1(R1610), .clock(clock), .in1(R1609));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1681 (.out1(R1682), .clock(clock), .in1(R1681));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1753 (.out1(R1754), .clock(clock), .in1(R1753));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1816 (.out1(R1817), .clock(clock), .in1(R1816));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1879 (.out1(R1880), .clock(clock), .in1(R1879));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1933 (.out1(R1934), .clock(clock), .in1(ifout126));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op1986 (.out1(R1987), .clock(clock), .in1(_111));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op129 (.out1(_112), .in1(C80_265_D), .in2(R1987));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op362 (.out1(R363), .clock(clock), .in1(R362));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op489 (.out1(R490), .clock(clock), .in1(R489));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op615 (.out1(R616), .clock(clock), .in1(R615));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op733 (.out1(R734), .clock(clock), .in1(R733));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op850 (.out1(R851), .clock(clock), .in1(R850));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op959 (.out1(R960), .clock(clock), .in1(R959));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1067 (.out1(R1068), .clock(clock), .in1(R1067));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1167 (.out1(R1168), .clock(clock), .in1(R1167));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1266 (.out1(R1267), .clock(clock), .in1(R1266));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1357 (.out1(R1358), .clock(clock), .in1(R1357));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1447 (.out1(R1448), .clock(clock), .in1(R1447));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1529 (.out1(R1530), .clock(clock), .in1(R1529));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1610 (.out1(R1611), .clock(clock), .in1(R1610));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1682 (.out1(R1683), .clock(clock), .in1(R1682));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1754 (.out1(R1755), .clock(clock), .in1(R1754));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1817 (.out1(R1818), .clock(clock), .in1(R1817));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1880 (.out1(R1881), .clock(clock), .in1(R1880));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1934 (.out1(R1935), .clock(clock), .in1(R1934));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op1987 (.out1(R1988), .clock(clock), .in1(_112));
  SRAM op130 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_113),.ADR(R1988));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op363 (.out1(R364), .clock(clock), .in1(R363));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op490 (.out1(R491), .clock(clock), .in1(R490));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op616 (.out1(R617), .clock(clock), .in1(R616));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op734 (.out1(R735), .clock(clock), .in1(R734));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op851 (.out1(R852), .clock(clock), .in1(R851));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op960 (.out1(R961), .clock(clock), .in1(R960));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1068 (.out1(R1069), .clock(clock), .in1(R1068));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1168 (.out1(R1169), .clock(clock), .in1(R1168));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1267 (.out1(R1268), .clock(clock), .in1(R1267));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1358 (.out1(R1359), .clock(clock), .in1(R1358));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1448 (.out1(R1449), .clock(clock), .in1(R1448));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1530 (.out1(R1531), .clock(clock), .in1(R1530));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1611 (.out1(R1612), .clock(clock), .in1(R1611));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1683 (.out1(R1684), .clock(clock), .in1(R1683));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1755 (.out1(R1756), .clock(clock), .in1(R1755));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1818 (.out1(R1819), .clock(clock), .in1(R1818));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1881 (.out1(R1882), .clock(clock), .in1(R1881));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1935 (.out1(R1936), .clock(clock), .in1(R1935));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1988 (.out1(R1989), .clock(clock), .in1(_113));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op131 (.out1(_114), .in1(R1989), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op364 (.out1(R365), .clock(clock), .in1(R364));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op491 (.out1(R492), .clock(clock), .in1(R491));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op617 (.out1(R618), .clock(clock), .in1(R617));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op735 (.out1(R736), .clock(clock), .in1(R735));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op852 (.out1(R853), .clock(clock), .in1(R852));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op961 (.out1(R962), .clock(clock), .in1(R961));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1069 (.out1(R1070), .clock(clock), .in1(R1069));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1169 (.out1(R1170), .clock(clock), .in1(R1169));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1268 (.out1(R1269), .clock(clock), .in1(R1268));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1359 (.out1(R1360), .clock(clock), .in1(R1359));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1449 (.out1(R1450), .clock(clock), .in1(R1449));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1531 (.out1(R1532), .clock(clock), .in1(R1531));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1612 (.out1(R1613), .clock(clock), .in1(R1612));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1684 (.out1(R1685), .clock(clock), .in1(R1684));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1756 (.out1(R1757), .clock(clock), .in1(R1756));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1819 (.out1(R1820), .clock(clock), .in1(R1819));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1882 (.out1(R1883), .clock(clock), .in1(R1882));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1936 (.out1(R1937), .clock(clock), .in1(R1936));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1989 (.out1(R1990), .clock(clock), .in1(_114));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(4), .BITSIZE_out1(32), .PRECISION(32)) op132 (.out1(_115), .in1(R1990), .in2(4 'd 8));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op365 (.out1(R366), .clock(clock), .in1(R365));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op492 (.out1(R493), .clock(clock), .in1(R492));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op618 (.out1(R619), .clock(clock), .in1(R618));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op736 (.out1(R737), .clock(clock), .in1(R736));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op853 (.out1(R854), .clock(clock), .in1(R853));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op962 (.out1(R963), .clock(clock), .in1(R962));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1070 (.out1(R1071), .clock(clock), .in1(R1070));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1170 (.out1(R1171), .clock(clock), .in1(R1170));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1269 (.out1(R1270), .clock(clock), .in1(R1269));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1360 (.out1(R1361), .clock(clock), .in1(R1360));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1450 (.out1(R1451), .clock(clock), .in1(R1450));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1532 (.out1(R1533), .clock(clock), .in1(R1532));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1613 (.out1(R1614), .clock(clock), .in1(R1613));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1685 (.out1(R1686), .clock(clock), .in1(R1685));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1757 (.out1(R1758), .clock(clock), .in1(R1757));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1820 (.out1(R1821), .clock(clock), .in1(R1820));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1883 (.out1(R1884), .clock(clock), .in1(R1883));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1937 (.out1(R1938), .clock(clock), .in1(R1937));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1990 (.out1(R1991), .clock(clock), .in1(_115));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op133 (.out1(_116), .in1(ip2_259_D), .in2(6 'd 40));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op134 (.out1(_117), .in1(_116));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(8), .BITSIZE_out1(32)) op135 (.out1(_118), .in1(_117), .in2(8 'd 255));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op136 (.out1(idx_268), .in1(R1991), .in2(_118));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op366 (.out1(R367), .clock(clock), .in1(R366));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op493 (.out1(R494), .clock(clock), .in1(R493));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op619 (.out1(R620), .clock(clock), .in1(R619));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op737 (.out1(R738), .clock(clock), .in1(R737));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op854 (.out1(R855), .clock(clock), .in1(R854));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op963 (.out1(R964), .clock(clock), .in1(R963));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1071 (.out1(R1072), .clock(clock), .in1(R1071));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1171 (.out1(R1172), .clock(clock), .in1(R1171));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1270 (.out1(R1271), .clock(clock), .in1(R1270));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1361 (.out1(R1362), .clock(clock), .in1(R1361));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1451 (.out1(R1452), .clock(clock), .in1(R1451));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1533 (.out1(R1534), .clock(clock), .in1(R1533));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1614 (.out1(R1615), .clock(clock), .in1(R1614));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1686 (.out1(R1687), .clock(clock), .in1(R1686));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1758 (.out1(R1759), .clock(clock), .in1(R1758));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1821 (.out1(R1822), .clock(clock), .in1(R1821));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1884 (.out1(R1885), .clock(clock), .in1(R1884));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1938 (.out1(R1939), .clock(clock), .in1(R1938));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1991 (.out1(R1992), .clock(clock), .in1(idx_268));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op137 (.out1(_119), .in1(R1992));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op138 (.out1(_120), .in1(_119), .in2(2 'd 2));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op367 (.out1(R368), .clock(clock), .in1(R367));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op494 (.out1(R495), .clock(clock), .in1(R494));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op620 (.out1(R621), .clock(clock), .in1(R620));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op738 (.out1(R739), .clock(clock), .in1(R738));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op855 (.out1(R856), .clock(clock), .in1(R855));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op964 (.out1(R965), .clock(clock), .in1(R964));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1072 (.out1(R1073), .clock(clock), .in1(R1072));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1172 (.out1(R1173), .clock(clock), .in1(R1172));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1271 (.out1(R1272), .clock(clock), .in1(R1271));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1362 (.out1(R1363), .clock(clock), .in1(R1362));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1452 (.out1(R1453), .clock(clock), .in1(R1452));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1534 (.out1(R1535), .clock(clock), .in1(R1534));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1615 (.out1(R1616), .clock(clock), .in1(R1615));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1687 (.out1(R1688), .clock(clock), .in1(R1687));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1759 (.out1(R1760), .clock(clock), .in1(R1759));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1822 (.out1(R1823), .clock(clock), .in1(R1822));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1885 (.out1(R1886), .clock(clock), .in1(R1885));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1939 (.out1(R1940), .clock(clock), .in1(R1939));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1992 (.out1(R1993), .clock(clock), .in1(R1992));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2037 (.out1(R2038), .clock(clock), .in1(_120));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op139 (.out1(_121), .in1(C88_269_D), .in2(R2038));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op368 (.out1(R369), .clock(clock), .in1(R368));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op495 (.out1(R496), .clock(clock), .in1(R495));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op621 (.out1(R622), .clock(clock), .in1(R621));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op739 (.out1(R740), .clock(clock), .in1(R739));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op856 (.out1(R857), .clock(clock), .in1(R856));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op965 (.out1(R966), .clock(clock), .in1(R965));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1073 (.out1(R1074), .clock(clock), .in1(R1073));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1173 (.out1(R1174), .clock(clock), .in1(R1173));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1272 (.out1(R1273), .clock(clock), .in1(R1272));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1363 (.out1(R1364), .clock(clock), .in1(R1363));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1453 (.out1(R1454), .clock(clock), .in1(R1453));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1535 (.out1(R1536), .clock(clock), .in1(R1535));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1616 (.out1(R1617), .clock(clock), .in1(R1616));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1688 (.out1(R1689), .clock(clock), .in1(R1688));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1760 (.out1(R1761), .clock(clock), .in1(R1760));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1823 (.out1(R1824), .clock(clock), .in1(R1823));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1886 (.out1(R1887), .clock(clock), .in1(R1886));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1940 (.out1(R1941), .clock(clock), .in1(R1940));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1993 (.out1(R1994), .clock(clock), .in1(R1993));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2038 (.out1(R2039), .clock(clock), .in1(_121));
  SRAM op140 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_122),.ADR(R2039));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op369 (.out1(R370), .clock(clock), .in1(R369));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op496 (.out1(R497), .clock(clock), .in1(R496));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op622 (.out1(R623), .clock(clock), .in1(R622));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op740 (.out1(R741), .clock(clock), .in1(R740));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op857 (.out1(R858), .clock(clock), .in1(R857));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op966 (.out1(R967), .clock(clock), .in1(R966));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1074 (.out1(R1075), .clock(clock), .in1(R1074));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1174 (.out1(R1175), .clock(clock), .in1(R1174));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1273 (.out1(R1274), .clock(clock), .in1(R1273));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1364 (.out1(R1365), .clock(clock), .in1(R1364));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1454 (.out1(R1455), .clock(clock), .in1(R1454));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1536 (.out1(R1537), .clock(clock), .in1(R1536));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1617 (.out1(R1618), .clock(clock), .in1(R1617));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1689 (.out1(R1690), .clock(clock), .in1(R1689));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1761 (.out1(R1762), .clock(clock), .in1(R1761));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1824 (.out1(R1825), .clock(clock), .in1(R1824));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1887 (.out1(R1888), .clock(clock), .in1(R1887));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1941 (.out1(R1942), .clock(clock), .in1(R1941));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1994 (.out1(R1995), .clock(clock), .in1(R1994));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2039 (.out1(R2040), .clock(clock), .in1(_122));
  NE_EXPR #(.BITSIZE_in1(32), .BITSIZE_in2(1),.BITSIZE_out1(1)) op141 (.out1(ifout141), .in1(R2040), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op142 (.out1(_123), .in1(R1995));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op143 (.out1(_124), .in1(_123), .in2(2 'd 2));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op370 (.out1(R371), .clock(clock), .in1(R370));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op497 (.out1(R498), .clock(clock), .in1(R497));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op623 (.out1(R624), .clock(clock), .in1(R623));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op741 (.out1(R742), .clock(clock), .in1(R741));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op858 (.out1(R859), .clock(clock), .in1(R858));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op967 (.out1(R968), .clock(clock), .in1(R967));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1075 (.out1(R1076), .clock(clock), .in1(R1075));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1175 (.out1(R1176), .clock(clock), .in1(R1175));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1274 (.out1(R1275), .clock(clock), .in1(R1274));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1365 (.out1(R1366), .clock(clock), .in1(R1365));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1455 (.out1(R1456), .clock(clock), .in1(R1455));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1537 (.out1(R1538), .clock(clock), .in1(R1537));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1618 (.out1(R1619), .clock(clock), .in1(R1618));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1690 (.out1(R1691), .clock(clock), .in1(R1690));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1762 (.out1(R1763), .clock(clock), .in1(R1762));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1825 (.out1(R1826), .clock(clock), .in1(R1825));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1888 (.out1(R1889), .clock(clock), .in1(R1888));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1942 (.out1(R1943), .clock(clock), .in1(R1942));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1995 (.out1(R1996), .clock(clock), .in1(R1995));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2040 (.out1(R2041), .clock(clock), .in1(ifout141));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2084 (.out1(R2085), .clock(clock), .in1(_124));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op144 (.out1(_125), .in1(C88_269_D), .in2(R2085));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op371 (.out1(R372), .clock(clock), .in1(R371));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op498 (.out1(R499), .clock(clock), .in1(R498));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op624 (.out1(R625), .clock(clock), .in1(R624));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op742 (.out1(R743), .clock(clock), .in1(R742));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op859 (.out1(R860), .clock(clock), .in1(R859));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op968 (.out1(R969), .clock(clock), .in1(R968));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1076 (.out1(R1077), .clock(clock), .in1(R1076));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1176 (.out1(R1177), .clock(clock), .in1(R1176));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1275 (.out1(R1276), .clock(clock), .in1(R1275));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1366 (.out1(R1367), .clock(clock), .in1(R1366));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1456 (.out1(R1457), .clock(clock), .in1(R1456));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1538 (.out1(R1539), .clock(clock), .in1(R1538));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1619 (.out1(R1620), .clock(clock), .in1(R1619));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1691 (.out1(R1692), .clock(clock), .in1(R1691));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1763 (.out1(R1764), .clock(clock), .in1(R1763));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1826 (.out1(R1827), .clock(clock), .in1(R1826));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1889 (.out1(R1890), .clock(clock), .in1(R1889));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1943 (.out1(R1944), .clock(clock), .in1(R1943));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1996 (.out1(R1997), .clock(clock), .in1(R1996));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2041 (.out1(R2042), .clock(clock), .in1(R2041));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2085 (.out1(R2086), .clock(clock), .in1(_125));
  SRAM op145 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_126),.ADR(R2086));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op372 (.out1(R373), .clock(clock), .in1(R372));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op499 (.out1(R500), .clock(clock), .in1(R499));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op625 (.out1(R626), .clock(clock), .in1(R625));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op743 (.out1(R744), .clock(clock), .in1(R743));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op860 (.out1(R861), .clock(clock), .in1(R860));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op969 (.out1(R970), .clock(clock), .in1(R969));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1077 (.out1(R1078), .clock(clock), .in1(R1077));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1177 (.out1(R1178), .clock(clock), .in1(R1177));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1276 (.out1(R1277), .clock(clock), .in1(R1276));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1367 (.out1(R1368), .clock(clock), .in1(R1367));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1457 (.out1(R1458), .clock(clock), .in1(R1457));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1539 (.out1(R1540), .clock(clock), .in1(R1539));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1620 (.out1(R1621), .clock(clock), .in1(R1620));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1692 (.out1(R1693), .clock(clock), .in1(R1692));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1764 (.out1(R1765), .clock(clock), .in1(R1764));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1827 (.out1(R1828), .clock(clock), .in1(R1827));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1890 (.out1(R1891), .clock(clock), .in1(R1890));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1944 (.out1(R1945), .clock(clock), .in1(R1944));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1997 (.out1(R1998), .clock(clock), .in1(R1997));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2042 (.out1(R2043), .clock(clock), .in1(R2042));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2086 (.out1(R2087), .clock(clock), .in1(_126));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op146 (.out1(_127), .in1(R2087), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op373 (.out1(R374), .clock(clock), .in1(R373));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op500 (.out1(R501), .clock(clock), .in1(R500));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op626 (.out1(R627), .clock(clock), .in1(R626));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op744 (.out1(R745), .clock(clock), .in1(R744));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op861 (.out1(R862), .clock(clock), .in1(R861));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op970 (.out1(R971), .clock(clock), .in1(R970));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1078 (.out1(R1079), .clock(clock), .in1(R1078));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1178 (.out1(R1179), .clock(clock), .in1(R1178));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1277 (.out1(R1278), .clock(clock), .in1(R1277));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1368 (.out1(R1369), .clock(clock), .in1(R1368));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1458 (.out1(R1459), .clock(clock), .in1(R1458));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1540 (.out1(R1541), .clock(clock), .in1(R1540));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1621 (.out1(R1622), .clock(clock), .in1(R1621));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1693 (.out1(R1694), .clock(clock), .in1(R1693));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1765 (.out1(R1766), .clock(clock), .in1(R1765));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1828 (.out1(R1829), .clock(clock), .in1(R1828));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1891 (.out1(R1892), .clock(clock), .in1(R1891));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1945 (.out1(R1946), .clock(clock), .in1(R1945));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1998 (.out1(R1999), .clock(clock), .in1(R1998));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2043 (.out1(R2044), .clock(clock), .in1(R2043));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2087 (.out1(R2088), .clock(clock), .in1(_127));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(4), .BITSIZE_out1(32), .PRECISION(32)) op147 (.out1(_128), .in1(R2088), .in2(4 'd 8));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op374 (.out1(R375), .clock(clock), .in1(R374));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op501 (.out1(R502), .clock(clock), .in1(R501));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op627 (.out1(R628), .clock(clock), .in1(R627));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op745 (.out1(R746), .clock(clock), .in1(R745));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op862 (.out1(R863), .clock(clock), .in1(R862));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op971 (.out1(R972), .clock(clock), .in1(R971));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1079 (.out1(R1080), .clock(clock), .in1(R1079));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1179 (.out1(R1180), .clock(clock), .in1(R1179));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1278 (.out1(R1279), .clock(clock), .in1(R1278));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1369 (.out1(R1370), .clock(clock), .in1(R1369));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1459 (.out1(R1460), .clock(clock), .in1(R1459));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1541 (.out1(R1542), .clock(clock), .in1(R1541));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1622 (.out1(R1623), .clock(clock), .in1(R1622));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1694 (.out1(R1695), .clock(clock), .in1(R1694));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1766 (.out1(R1767), .clock(clock), .in1(R1766));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1829 (.out1(R1830), .clock(clock), .in1(R1829));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1892 (.out1(R1893), .clock(clock), .in1(R1892));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1946 (.out1(R1947), .clock(clock), .in1(R1946));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1999 (.out1(R2000), .clock(clock), .in1(R1999));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2044 (.out1(R2045), .clock(clock), .in1(R2044));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2088 (.out1(R2089), .clock(clock), .in1(_128));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op148 (.out1(_129), .in1(ip2_259_D), .in2(6 'd 32));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op149 (.out1(_130), .in1(_129));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(8), .BITSIZE_out1(32)) op150 (.out1(_131), .in1(_130), .in2(8 'd 255));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op151 (.out1(idx_272), .in1(R2089), .in2(_131));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op375 (.out1(R376), .clock(clock), .in1(R375));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op502 (.out1(R503), .clock(clock), .in1(R502));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op628 (.out1(R629), .clock(clock), .in1(R628));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op746 (.out1(R747), .clock(clock), .in1(R746));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op863 (.out1(R864), .clock(clock), .in1(R863));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op972 (.out1(R973), .clock(clock), .in1(R972));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1080 (.out1(R1081), .clock(clock), .in1(R1080));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1180 (.out1(R1181), .clock(clock), .in1(R1180));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1279 (.out1(R1280), .clock(clock), .in1(R1279));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1370 (.out1(R1371), .clock(clock), .in1(R1370));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1460 (.out1(R1461), .clock(clock), .in1(R1460));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1542 (.out1(R1543), .clock(clock), .in1(R1542));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1623 (.out1(R1624), .clock(clock), .in1(R1623));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1695 (.out1(R1696), .clock(clock), .in1(R1695));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1767 (.out1(R1768), .clock(clock), .in1(R1767));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1830 (.out1(R1831), .clock(clock), .in1(R1830));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1893 (.out1(R1894), .clock(clock), .in1(R1893));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1947 (.out1(R1948), .clock(clock), .in1(R1947));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2000 (.out1(R2001), .clock(clock), .in1(R2000));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2045 (.out1(R2046), .clock(clock), .in1(R2045));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2089 (.out1(R2090), .clock(clock), .in1(idx_272));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op152 (.out1(_132), .in1(R2090));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op153 (.out1(_133), .in1(_132), .in2(2 'd 2));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op376 (.out1(R377), .clock(clock), .in1(R376));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op503 (.out1(R504), .clock(clock), .in1(R503));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op629 (.out1(R630), .clock(clock), .in1(R629));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op747 (.out1(R748), .clock(clock), .in1(R747));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op864 (.out1(R865), .clock(clock), .in1(R864));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op973 (.out1(R974), .clock(clock), .in1(R973));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1081 (.out1(R1082), .clock(clock), .in1(R1081));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1181 (.out1(R1182), .clock(clock), .in1(R1181));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1280 (.out1(R1281), .clock(clock), .in1(R1280));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1371 (.out1(R1372), .clock(clock), .in1(R1371));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1461 (.out1(R1462), .clock(clock), .in1(R1461));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1543 (.out1(R1544), .clock(clock), .in1(R1543));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1624 (.out1(R1625), .clock(clock), .in1(R1624));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1696 (.out1(R1697), .clock(clock), .in1(R1696));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1768 (.out1(R1769), .clock(clock), .in1(R1768));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1831 (.out1(R1832), .clock(clock), .in1(R1831));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1894 (.out1(R1895), .clock(clock), .in1(R1894));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1948 (.out1(R1949), .clock(clock), .in1(R1948));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2001 (.out1(R2002), .clock(clock), .in1(R2001));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2046 (.out1(R2047), .clock(clock), .in1(R2046));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2090 (.out1(R2091), .clock(clock), .in1(R2090));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2126 (.out1(R2127), .clock(clock), .in1(_133));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op154 (.out1(_134), .in1(C96_273_D), .in2(R2127));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op377 (.out1(R378), .clock(clock), .in1(R377));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op504 (.out1(R505), .clock(clock), .in1(R504));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op630 (.out1(R631), .clock(clock), .in1(R630));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op748 (.out1(R749), .clock(clock), .in1(R748));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op865 (.out1(R866), .clock(clock), .in1(R865));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op974 (.out1(R975), .clock(clock), .in1(R974));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1082 (.out1(R1083), .clock(clock), .in1(R1082));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1182 (.out1(R1183), .clock(clock), .in1(R1182));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1281 (.out1(R1282), .clock(clock), .in1(R1281));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1372 (.out1(R1373), .clock(clock), .in1(R1372));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1462 (.out1(R1463), .clock(clock), .in1(R1462));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1544 (.out1(R1545), .clock(clock), .in1(R1544));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1625 (.out1(R1626), .clock(clock), .in1(R1625));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1697 (.out1(R1698), .clock(clock), .in1(R1697));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1769 (.out1(R1770), .clock(clock), .in1(R1769));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1832 (.out1(R1833), .clock(clock), .in1(R1832));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1895 (.out1(R1896), .clock(clock), .in1(R1895));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1949 (.out1(R1950), .clock(clock), .in1(R1949));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2002 (.out1(R2003), .clock(clock), .in1(R2002));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2047 (.out1(R2048), .clock(clock), .in1(R2047));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2091 (.out1(R2092), .clock(clock), .in1(R2091));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2127 (.out1(R2128), .clock(clock), .in1(_134));
  SRAM op155 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_135),.ADR(R2128));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op378 (.out1(R379), .clock(clock), .in1(R378));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op505 (.out1(R506), .clock(clock), .in1(R505));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op631 (.out1(R632), .clock(clock), .in1(R631));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op749 (.out1(R750), .clock(clock), .in1(R749));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op866 (.out1(R867), .clock(clock), .in1(R866));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op975 (.out1(R976), .clock(clock), .in1(R975));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1083 (.out1(R1084), .clock(clock), .in1(R1083));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1183 (.out1(R1184), .clock(clock), .in1(R1183));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1282 (.out1(R1283), .clock(clock), .in1(R1282));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1373 (.out1(R1374), .clock(clock), .in1(R1373));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1463 (.out1(R1464), .clock(clock), .in1(R1463));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1545 (.out1(R1546), .clock(clock), .in1(R1545));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1626 (.out1(R1627), .clock(clock), .in1(R1626));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1698 (.out1(R1699), .clock(clock), .in1(R1698));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1770 (.out1(R1771), .clock(clock), .in1(R1770));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1833 (.out1(R1834), .clock(clock), .in1(R1833));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1896 (.out1(R1897), .clock(clock), .in1(R1896));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1950 (.out1(R1951), .clock(clock), .in1(R1950));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2003 (.out1(R2004), .clock(clock), .in1(R2003));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2048 (.out1(R2049), .clock(clock), .in1(R2048));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2092 (.out1(R2093), .clock(clock), .in1(R2092));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2128 (.out1(R2129), .clock(clock), .in1(_135));
  NE_EXPR #(.BITSIZE_in1(32), .BITSIZE_in2(1),.BITSIZE_out1(1)) op156 (.out1(ifout156), .in1(R2129), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op157 (.out1(_136), .in1(R2093));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op158 (.out1(_137), .in1(_136), .in2(2 'd 2));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op379 (.out1(R380), .clock(clock), .in1(R379));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op506 (.out1(R507), .clock(clock), .in1(R506));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op632 (.out1(R633), .clock(clock), .in1(R632));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op750 (.out1(R751), .clock(clock), .in1(R750));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op867 (.out1(R868), .clock(clock), .in1(R867));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op976 (.out1(R977), .clock(clock), .in1(R976));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1084 (.out1(R1085), .clock(clock), .in1(R1084));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1184 (.out1(R1185), .clock(clock), .in1(R1184));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1283 (.out1(R1284), .clock(clock), .in1(R1283));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1374 (.out1(R1375), .clock(clock), .in1(R1374));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1464 (.out1(R1465), .clock(clock), .in1(R1464));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1546 (.out1(R1547), .clock(clock), .in1(R1546));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1627 (.out1(R1628), .clock(clock), .in1(R1627));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1699 (.out1(R1700), .clock(clock), .in1(R1699));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1771 (.out1(R1772), .clock(clock), .in1(R1771));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1834 (.out1(R1835), .clock(clock), .in1(R1834));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1897 (.out1(R1898), .clock(clock), .in1(R1897));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1951 (.out1(R1952), .clock(clock), .in1(R1951));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2004 (.out1(R2005), .clock(clock), .in1(R2004));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2049 (.out1(R2050), .clock(clock), .in1(R2049));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2093 (.out1(R2094), .clock(clock), .in1(R2093));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2129 (.out1(R2130), .clock(clock), .in1(ifout156));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2164 (.out1(R2165), .clock(clock), .in1(_137));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op159 (.out1(_138), .in1(C96_273_D), .in2(R2165));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op380 (.out1(R381), .clock(clock), .in1(R380));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op507 (.out1(R508), .clock(clock), .in1(R507));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op633 (.out1(R634), .clock(clock), .in1(R633));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op751 (.out1(R752), .clock(clock), .in1(R751));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op868 (.out1(R869), .clock(clock), .in1(R868));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op977 (.out1(R978), .clock(clock), .in1(R977));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1085 (.out1(R1086), .clock(clock), .in1(R1085));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1185 (.out1(R1186), .clock(clock), .in1(R1185));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1284 (.out1(R1285), .clock(clock), .in1(R1284));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1375 (.out1(R1376), .clock(clock), .in1(R1375));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1465 (.out1(R1466), .clock(clock), .in1(R1465));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1547 (.out1(R1548), .clock(clock), .in1(R1547));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1628 (.out1(R1629), .clock(clock), .in1(R1628));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1700 (.out1(R1701), .clock(clock), .in1(R1700));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1772 (.out1(R1773), .clock(clock), .in1(R1772));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1835 (.out1(R1836), .clock(clock), .in1(R1835));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1898 (.out1(R1899), .clock(clock), .in1(R1898));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1952 (.out1(R1953), .clock(clock), .in1(R1952));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2005 (.out1(R2006), .clock(clock), .in1(R2005));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2050 (.out1(R2051), .clock(clock), .in1(R2050));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2094 (.out1(R2095), .clock(clock), .in1(R2094));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2130 (.out1(R2131), .clock(clock), .in1(R2130));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2165 (.out1(R2166), .clock(clock), .in1(_138));
  SRAM op160 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_139),.ADR(R2166));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op381 (.out1(R382), .clock(clock), .in1(R381));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op508 (.out1(R509), .clock(clock), .in1(R508));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op634 (.out1(R635), .clock(clock), .in1(R634));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op752 (.out1(R753), .clock(clock), .in1(R752));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op869 (.out1(R870), .clock(clock), .in1(R869));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op978 (.out1(R979), .clock(clock), .in1(R978));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1086 (.out1(R1087), .clock(clock), .in1(R1086));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1186 (.out1(R1187), .clock(clock), .in1(R1186));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1285 (.out1(R1286), .clock(clock), .in1(R1285));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1376 (.out1(R1377), .clock(clock), .in1(R1376));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1466 (.out1(R1467), .clock(clock), .in1(R1466));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1548 (.out1(R1549), .clock(clock), .in1(R1548));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1629 (.out1(R1630), .clock(clock), .in1(R1629));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1701 (.out1(R1702), .clock(clock), .in1(R1701));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1773 (.out1(R1774), .clock(clock), .in1(R1773));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1836 (.out1(R1837), .clock(clock), .in1(R1836));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1899 (.out1(R1900), .clock(clock), .in1(R1899));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1953 (.out1(R1954), .clock(clock), .in1(R1953));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2006 (.out1(R2007), .clock(clock), .in1(R2006));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2051 (.out1(R2052), .clock(clock), .in1(R2051));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2095 (.out1(R2096), .clock(clock), .in1(R2095));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2131 (.out1(R2132), .clock(clock), .in1(R2131));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2166 (.out1(R2167), .clock(clock), .in1(_139));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op161 (.out1(_140), .in1(R2167), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op382 (.out1(R383), .clock(clock), .in1(R382));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op509 (.out1(R510), .clock(clock), .in1(R509));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op635 (.out1(R636), .clock(clock), .in1(R635));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op753 (.out1(R754), .clock(clock), .in1(R753));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op870 (.out1(R871), .clock(clock), .in1(R870));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op979 (.out1(R980), .clock(clock), .in1(R979));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1087 (.out1(R1088), .clock(clock), .in1(R1087));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1187 (.out1(R1188), .clock(clock), .in1(R1187));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1286 (.out1(R1287), .clock(clock), .in1(R1286));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1377 (.out1(R1378), .clock(clock), .in1(R1377));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1467 (.out1(R1468), .clock(clock), .in1(R1467));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1549 (.out1(R1550), .clock(clock), .in1(R1549));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1630 (.out1(R1631), .clock(clock), .in1(R1630));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1702 (.out1(R1703), .clock(clock), .in1(R1702));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1774 (.out1(R1775), .clock(clock), .in1(R1774));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1837 (.out1(R1838), .clock(clock), .in1(R1837));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1900 (.out1(R1901), .clock(clock), .in1(R1900));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1954 (.out1(R1955), .clock(clock), .in1(R1954));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2007 (.out1(R2008), .clock(clock), .in1(R2007));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2052 (.out1(R2053), .clock(clock), .in1(R2052));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2096 (.out1(R2097), .clock(clock), .in1(R2096));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2132 (.out1(R2133), .clock(clock), .in1(R2132));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2167 (.out1(R2168), .clock(clock), .in1(_140));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(4), .BITSIZE_out1(32), .PRECISION(32)) op162 (.out1(_141), .in1(R2168), .in2(4 'd 8));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op383 (.out1(R384), .clock(clock), .in1(R383));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op510 (.out1(R511), .clock(clock), .in1(R510));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op636 (.out1(R637), .clock(clock), .in1(R636));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op754 (.out1(R755), .clock(clock), .in1(R754));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op871 (.out1(R872), .clock(clock), .in1(R871));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op980 (.out1(R981), .clock(clock), .in1(R980));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1088 (.out1(R1089), .clock(clock), .in1(R1088));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1188 (.out1(R1189), .clock(clock), .in1(R1188));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1287 (.out1(R1288), .clock(clock), .in1(R1287));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1378 (.out1(R1379), .clock(clock), .in1(R1378));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1468 (.out1(R1469), .clock(clock), .in1(R1468));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1550 (.out1(R1551), .clock(clock), .in1(R1550));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1631 (.out1(R1632), .clock(clock), .in1(R1631));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1703 (.out1(R1704), .clock(clock), .in1(R1703));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1775 (.out1(R1776), .clock(clock), .in1(R1775));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1838 (.out1(R1839), .clock(clock), .in1(R1838));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1901 (.out1(R1902), .clock(clock), .in1(R1901));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1955 (.out1(R1956), .clock(clock), .in1(R1955));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2008 (.out1(R2009), .clock(clock), .in1(R2008));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2053 (.out1(R2054), .clock(clock), .in1(R2053));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2097 (.out1(R2098), .clock(clock), .in1(R2097));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2133 (.out1(R2134), .clock(clock), .in1(R2133));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2168 (.out1(R2169), .clock(clock), .in1(_141));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(5), .BITSIZE_out1(64), .PRECISION(64)) op163 (.out1(_142), .in1(ip2_259_D), .in2(5 'd 24));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op164 (.out1(_143), .in1(_142));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(8), .BITSIZE_out1(32)) op165 (.out1(_144), .in1(_143), .in2(8 'd 255));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op166 (.out1(idx_276), .in1(R2169), .in2(_144));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op384 (.out1(R385), .clock(clock), .in1(R384));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op511 (.out1(R512), .clock(clock), .in1(R511));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op637 (.out1(R638), .clock(clock), .in1(R637));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op755 (.out1(R756), .clock(clock), .in1(R755));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op872 (.out1(R873), .clock(clock), .in1(R872));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op981 (.out1(R982), .clock(clock), .in1(R981));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1089 (.out1(R1090), .clock(clock), .in1(R1089));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1189 (.out1(R1190), .clock(clock), .in1(R1189));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1288 (.out1(R1289), .clock(clock), .in1(R1288));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1379 (.out1(R1380), .clock(clock), .in1(R1379));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1469 (.out1(R1470), .clock(clock), .in1(R1469));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1551 (.out1(R1552), .clock(clock), .in1(R1551));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1632 (.out1(R1633), .clock(clock), .in1(R1632));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1704 (.out1(R1705), .clock(clock), .in1(R1704));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1776 (.out1(R1777), .clock(clock), .in1(R1776));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1839 (.out1(R1840), .clock(clock), .in1(R1839));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1902 (.out1(R1903), .clock(clock), .in1(R1902));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1956 (.out1(R1957), .clock(clock), .in1(R1956));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2009 (.out1(R2010), .clock(clock), .in1(R2009));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2054 (.out1(R2055), .clock(clock), .in1(R2054));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2098 (.out1(R2099), .clock(clock), .in1(R2098));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2134 (.out1(R2135), .clock(clock), .in1(R2134));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2169 (.out1(R2170), .clock(clock), .in1(idx_276));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op167 (.out1(_145), .in1(R2170));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op168 (.out1(_146), .in1(_145), .in2(2 'd 2));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op385 (.out1(R386), .clock(clock), .in1(R385));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op512 (.out1(R513), .clock(clock), .in1(R512));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op638 (.out1(R639), .clock(clock), .in1(R638));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op756 (.out1(R757), .clock(clock), .in1(R756));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op873 (.out1(R874), .clock(clock), .in1(R873));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op982 (.out1(R983), .clock(clock), .in1(R982));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1090 (.out1(R1091), .clock(clock), .in1(R1090));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1190 (.out1(R1191), .clock(clock), .in1(R1190));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1289 (.out1(R1290), .clock(clock), .in1(R1289));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1380 (.out1(R1381), .clock(clock), .in1(R1380));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1470 (.out1(R1471), .clock(clock), .in1(R1470));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1552 (.out1(R1553), .clock(clock), .in1(R1552));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1633 (.out1(R1634), .clock(clock), .in1(R1633));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1705 (.out1(R1706), .clock(clock), .in1(R1705));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1777 (.out1(R1778), .clock(clock), .in1(R1777));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1840 (.out1(R1841), .clock(clock), .in1(R1840));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1903 (.out1(R1904), .clock(clock), .in1(R1903));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1957 (.out1(R1958), .clock(clock), .in1(R1957));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2010 (.out1(R2011), .clock(clock), .in1(R2010));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2055 (.out1(R2056), .clock(clock), .in1(R2055));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2099 (.out1(R2100), .clock(clock), .in1(R2099));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2135 (.out1(R2136), .clock(clock), .in1(R2135));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2170 (.out1(R2171), .clock(clock), .in1(R2170));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2197 (.out1(R2198), .clock(clock), .in1(_146));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op169 (.out1(_147), .in1(C104_277_D), .in2(R2198));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op386 (.out1(R387), .clock(clock), .in1(R386));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op513 (.out1(R514), .clock(clock), .in1(R513));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op639 (.out1(R640), .clock(clock), .in1(R639));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op757 (.out1(R758), .clock(clock), .in1(R757));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op874 (.out1(R875), .clock(clock), .in1(R874));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op983 (.out1(R984), .clock(clock), .in1(R983));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1091 (.out1(R1092), .clock(clock), .in1(R1091));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1191 (.out1(R1192), .clock(clock), .in1(R1191));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1290 (.out1(R1291), .clock(clock), .in1(R1290));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1381 (.out1(R1382), .clock(clock), .in1(R1381));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1471 (.out1(R1472), .clock(clock), .in1(R1471));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1553 (.out1(R1554), .clock(clock), .in1(R1553));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1634 (.out1(R1635), .clock(clock), .in1(R1634));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1706 (.out1(R1707), .clock(clock), .in1(R1706));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1778 (.out1(R1779), .clock(clock), .in1(R1778));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1841 (.out1(R1842), .clock(clock), .in1(R1841));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1904 (.out1(R1905), .clock(clock), .in1(R1904));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1958 (.out1(R1959), .clock(clock), .in1(R1958));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2011 (.out1(R2012), .clock(clock), .in1(R2011));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2056 (.out1(R2057), .clock(clock), .in1(R2056));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2100 (.out1(R2101), .clock(clock), .in1(R2100));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2136 (.out1(R2137), .clock(clock), .in1(R2136));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2171 (.out1(R2172), .clock(clock), .in1(R2171));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2198 (.out1(R2199), .clock(clock), .in1(_147));
  SRAM op170 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_148),.ADR(R2199));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op387 (.out1(R388), .clock(clock), .in1(R387));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op514 (.out1(R515), .clock(clock), .in1(R514));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op640 (.out1(R641), .clock(clock), .in1(R640));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op758 (.out1(R759), .clock(clock), .in1(R758));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op875 (.out1(R876), .clock(clock), .in1(R875));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op984 (.out1(R985), .clock(clock), .in1(R984));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1092 (.out1(R1093), .clock(clock), .in1(R1092));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1192 (.out1(R1193), .clock(clock), .in1(R1192));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1291 (.out1(R1292), .clock(clock), .in1(R1291));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1382 (.out1(R1383), .clock(clock), .in1(R1382));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1472 (.out1(R1473), .clock(clock), .in1(R1472));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1554 (.out1(R1555), .clock(clock), .in1(R1554));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1635 (.out1(R1636), .clock(clock), .in1(R1635));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1707 (.out1(R1708), .clock(clock), .in1(R1707));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1779 (.out1(R1780), .clock(clock), .in1(R1779));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1842 (.out1(R1843), .clock(clock), .in1(R1842));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1905 (.out1(R1906), .clock(clock), .in1(R1905));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1959 (.out1(R1960), .clock(clock), .in1(R1959));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2012 (.out1(R2013), .clock(clock), .in1(R2012));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2057 (.out1(R2058), .clock(clock), .in1(R2057));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2101 (.out1(R2102), .clock(clock), .in1(R2101));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2137 (.out1(R2138), .clock(clock), .in1(R2137));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2172 (.out1(R2173), .clock(clock), .in1(R2172));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2199 (.out1(R2200), .clock(clock), .in1(_148));
  NE_EXPR #(.BITSIZE_in1(32), .BITSIZE_in2(1),.BITSIZE_out1(1)) op171 (.out1(ifout171), .in1(R2200), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op172 (.out1(_149), .in1(R2173));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op173 (.out1(_150), .in1(_149), .in2(2 'd 2));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op388 (.out1(R389), .clock(clock), .in1(R388));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op515 (.out1(R516), .clock(clock), .in1(R515));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op641 (.out1(R642), .clock(clock), .in1(R641));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op759 (.out1(R760), .clock(clock), .in1(R759));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op876 (.out1(R877), .clock(clock), .in1(R876));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op985 (.out1(R986), .clock(clock), .in1(R985));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1093 (.out1(R1094), .clock(clock), .in1(R1093));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1193 (.out1(R1194), .clock(clock), .in1(R1193));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1292 (.out1(R1293), .clock(clock), .in1(R1292));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1383 (.out1(R1384), .clock(clock), .in1(R1383));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1473 (.out1(R1474), .clock(clock), .in1(R1473));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1555 (.out1(R1556), .clock(clock), .in1(R1555));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1636 (.out1(R1637), .clock(clock), .in1(R1636));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1708 (.out1(R1709), .clock(clock), .in1(R1708));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1780 (.out1(R1781), .clock(clock), .in1(R1780));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1843 (.out1(R1844), .clock(clock), .in1(R1843));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1906 (.out1(R1907), .clock(clock), .in1(R1906));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1960 (.out1(R1961), .clock(clock), .in1(R1960));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2013 (.out1(R2014), .clock(clock), .in1(R2013));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2058 (.out1(R2059), .clock(clock), .in1(R2058));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2102 (.out1(R2103), .clock(clock), .in1(R2102));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2138 (.out1(R2139), .clock(clock), .in1(R2138));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2173 (.out1(R2174), .clock(clock), .in1(R2173));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2200 (.out1(R2201), .clock(clock), .in1(ifout171));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2226 (.out1(R2227), .clock(clock), .in1(_150));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op174 (.out1(_151), .in1(C104_277_D), .in2(R2227));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op389 (.out1(R390), .clock(clock), .in1(R389));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op516 (.out1(R517), .clock(clock), .in1(R516));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op642 (.out1(R643), .clock(clock), .in1(R642));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op760 (.out1(R761), .clock(clock), .in1(R760));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op877 (.out1(R878), .clock(clock), .in1(R877));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op986 (.out1(R987), .clock(clock), .in1(R986));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1094 (.out1(R1095), .clock(clock), .in1(R1094));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1194 (.out1(R1195), .clock(clock), .in1(R1194));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1293 (.out1(R1294), .clock(clock), .in1(R1293));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1384 (.out1(R1385), .clock(clock), .in1(R1384));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1474 (.out1(R1475), .clock(clock), .in1(R1474));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1556 (.out1(R1557), .clock(clock), .in1(R1556));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1637 (.out1(R1638), .clock(clock), .in1(R1637));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1709 (.out1(R1710), .clock(clock), .in1(R1709));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1781 (.out1(R1782), .clock(clock), .in1(R1781));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1844 (.out1(R1845), .clock(clock), .in1(R1844));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1907 (.out1(R1908), .clock(clock), .in1(R1907));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1961 (.out1(R1962), .clock(clock), .in1(R1961));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2014 (.out1(R2015), .clock(clock), .in1(R2014));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2059 (.out1(R2060), .clock(clock), .in1(R2059));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2103 (.out1(R2104), .clock(clock), .in1(R2103));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2139 (.out1(R2140), .clock(clock), .in1(R2139));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2174 (.out1(R2175), .clock(clock), .in1(R2174));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2201 (.out1(R2202), .clock(clock), .in1(R2201));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2227 (.out1(R2228), .clock(clock), .in1(_151));
  SRAM op175 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_152),.ADR(R2228));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op390 (.out1(R391), .clock(clock), .in1(R390));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op517 (.out1(R518), .clock(clock), .in1(R517));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op643 (.out1(R644), .clock(clock), .in1(R643));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op761 (.out1(R762), .clock(clock), .in1(R761));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op878 (.out1(R879), .clock(clock), .in1(R878));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op987 (.out1(R988), .clock(clock), .in1(R987));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1095 (.out1(R1096), .clock(clock), .in1(R1095));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1195 (.out1(R1196), .clock(clock), .in1(R1195));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1294 (.out1(R1295), .clock(clock), .in1(R1294));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1385 (.out1(R1386), .clock(clock), .in1(R1385));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1475 (.out1(R1476), .clock(clock), .in1(R1475));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1557 (.out1(R1558), .clock(clock), .in1(R1557));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1638 (.out1(R1639), .clock(clock), .in1(R1638));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1710 (.out1(R1711), .clock(clock), .in1(R1710));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1782 (.out1(R1783), .clock(clock), .in1(R1782));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1845 (.out1(R1846), .clock(clock), .in1(R1845));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1908 (.out1(R1909), .clock(clock), .in1(R1908));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1962 (.out1(R1963), .clock(clock), .in1(R1962));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2015 (.out1(R2016), .clock(clock), .in1(R2015));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2060 (.out1(R2061), .clock(clock), .in1(R2060));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2104 (.out1(R2105), .clock(clock), .in1(R2104));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2140 (.out1(R2141), .clock(clock), .in1(R2140));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2175 (.out1(R2176), .clock(clock), .in1(R2175));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2202 (.out1(R2203), .clock(clock), .in1(R2202));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2228 (.out1(R2229), .clock(clock), .in1(_152));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op176 (.out1(_153), .in1(R2229), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op391 (.out1(R392), .clock(clock), .in1(R391));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op518 (.out1(R519), .clock(clock), .in1(R518));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op644 (.out1(R645), .clock(clock), .in1(R644));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op762 (.out1(R763), .clock(clock), .in1(R762));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op879 (.out1(R880), .clock(clock), .in1(R879));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op988 (.out1(R989), .clock(clock), .in1(R988));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1096 (.out1(R1097), .clock(clock), .in1(R1096));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1196 (.out1(R1197), .clock(clock), .in1(R1196));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1295 (.out1(R1296), .clock(clock), .in1(R1295));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1386 (.out1(R1387), .clock(clock), .in1(R1386));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1476 (.out1(R1477), .clock(clock), .in1(R1476));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1558 (.out1(R1559), .clock(clock), .in1(R1558));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1639 (.out1(R1640), .clock(clock), .in1(R1639));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1711 (.out1(R1712), .clock(clock), .in1(R1711));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1783 (.out1(R1784), .clock(clock), .in1(R1783));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1846 (.out1(R1847), .clock(clock), .in1(R1846));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1909 (.out1(R1910), .clock(clock), .in1(R1909));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1963 (.out1(R1964), .clock(clock), .in1(R1963));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2016 (.out1(R2017), .clock(clock), .in1(R2016));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2061 (.out1(R2062), .clock(clock), .in1(R2061));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2105 (.out1(R2106), .clock(clock), .in1(R2105));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2141 (.out1(R2142), .clock(clock), .in1(R2141));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2176 (.out1(R2177), .clock(clock), .in1(R2176));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2203 (.out1(R2204), .clock(clock), .in1(R2203));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2229 (.out1(R2230), .clock(clock), .in1(_153));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(4), .BITSIZE_out1(32), .PRECISION(32)) op177 (.out1(_154), .in1(R2230), .in2(4 'd 8));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op392 (.out1(R393), .clock(clock), .in1(R392));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op519 (.out1(R520), .clock(clock), .in1(R519));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op645 (.out1(R646), .clock(clock), .in1(R645));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op763 (.out1(R764), .clock(clock), .in1(R763));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op880 (.out1(R881), .clock(clock), .in1(R880));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op989 (.out1(R990), .clock(clock), .in1(R989));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1097 (.out1(R1098), .clock(clock), .in1(R1097));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1197 (.out1(R1198), .clock(clock), .in1(R1197));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1296 (.out1(R1297), .clock(clock), .in1(R1296));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1387 (.out1(R1388), .clock(clock), .in1(R1387));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1477 (.out1(R1478), .clock(clock), .in1(R1477));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1559 (.out1(R1560), .clock(clock), .in1(R1559));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1640 (.out1(R1641), .clock(clock), .in1(R1640));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1712 (.out1(R1713), .clock(clock), .in1(R1712));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1784 (.out1(R1785), .clock(clock), .in1(R1784));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1847 (.out1(R1848), .clock(clock), .in1(R1847));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1910 (.out1(R1911), .clock(clock), .in1(R1910));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1964 (.out1(R1965), .clock(clock), .in1(R1964));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2017 (.out1(R2018), .clock(clock), .in1(R2017));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2062 (.out1(R2063), .clock(clock), .in1(R2062));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2106 (.out1(R2107), .clock(clock), .in1(R2106));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2142 (.out1(R2143), .clock(clock), .in1(R2142));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2177 (.out1(R2178), .clock(clock), .in1(R2177));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2204 (.out1(R2205), .clock(clock), .in1(R2204));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2230 (.out1(R2231), .clock(clock), .in1(_154));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(5), .BITSIZE_out1(64), .PRECISION(64)) op178 (.out1(_155), .in1(ip2_259_D), .in2(5 'd 16));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op179 (.out1(_156), .in1(_155));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(8), .BITSIZE_out1(32)) op180 (.out1(_157), .in1(_156), .in2(8 'd 255));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op181 (.out1(idx_280), .in1(R2231), .in2(_157));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op393 (.out1(R394), .clock(clock), .in1(R393));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op520 (.out1(R521), .clock(clock), .in1(R520));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op646 (.out1(R647), .clock(clock), .in1(R646));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op764 (.out1(R765), .clock(clock), .in1(R764));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op881 (.out1(R882), .clock(clock), .in1(R881));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op990 (.out1(R991), .clock(clock), .in1(R990));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1098 (.out1(R1099), .clock(clock), .in1(R1098));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1198 (.out1(R1199), .clock(clock), .in1(R1198));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1297 (.out1(R1298), .clock(clock), .in1(R1297));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1388 (.out1(R1389), .clock(clock), .in1(R1388));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1478 (.out1(R1479), .clock(clock), .in1(R1478));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1560 (.out1(R1561), .clock(clock), .in1(R1560));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1641 (.out1(R1642), .clock(clock), .in1(R1641));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1713 (.out1(R1714), .clock(clock), .in1(R1713));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1785 (.out1(R1786), .clock(clock), .in1(R1785));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1848 (.out1(R1849), .clock(clock), .in1(R1848));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1911 (.out1(R1912), .clock(clock), .in1(R1911));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1965 (.out1(R1966), .clock(clock), .in1(R1965));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2018 (.out1(R2019), .clock(clock), .in1(R2018));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2063 (.out1(R2064), .clock(clock), .in1(R2063));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2107 (.out1(R2108), .clock(clock), .in1(R2107));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2143 (.out1(R2144), .clock(clock), .in1(R2143));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2178 (.out1(R2179), .clock(clock), .in1(R2178));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2205 (.out1(R2206), .clock(clock), .in1(R2205));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2231 (.out1(R2232), .clock(clock), .in1(idx_280));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op182 (.out1(_158), .in1(R2232));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op183 (.out1(_159), .in1(_158), .in2(2 'd 2));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op394 (.out1(R395), .clock(clock), .in1(R394));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op521 (.out1(R522), .clock(clock), .in1(R521));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op647 (.out1(R648), .clock(clock), .in1(R647));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op765 (.out1(R766), .clock(clock), .in1(R765));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op882 (.out1(R883), .clock(clock), .in1(R882));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op991 (.out1(R992), .clock(clock), .in1(R991));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1099 (.out1(R1100), .clock(clock), .in1(R1099));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1199 (.out1(R1200), .clock(clock), .in1(R1199));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1298 (.out1(R1299), .clock(clock), .in1(R1298));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1389 (.out1(R1390), .clock(clock), .in1(R1389));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1479 (.out1(R1480), .clock(clock), .in1(R1479));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1561 (.out1(R1562), .clock(clock), .in1(R1561));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1642 (.out1(R1643), .clock(clock), .in1(R1642));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1714 (.out1(R1715), .clock(clock), .in1(R1714));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1786 (.out1(R1787), .clock(clock), .in1(R1786));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1849 (.out1(R1850), .clock(clock), .in1(R1849));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1912 (.out1(R1913), .clock(clock), .in1(R1912));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1966 (.out1(R1967), .clock(clock), .in1(R1966));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2019 (.out1(R2020), .clock(clock), .in1(R2019));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2064 (.out1(R2065), .clock(clock), .in1(R2064));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2108 (.out1(R2109), .clock(clock), .in1(R2108));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2144 (.out1(R2145), .clock(clock), .in1(R2144));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2179 (.out1(R2180), .clock(clock), .in1(R2179));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2206 (.out1(R2207), .clock(clock), .in1(R2206));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2232 (.out1(R2233), .clock(clock), .in1(R2232));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2250 (.out1(R2251), .clock(clock), .in1(_159));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op184 (.out1(_160), .in1(C112_281_D), .in2(R2251));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op395 (.out1(R396), .clock(clock), .in1(R395));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op522 (.out1(R523), .clock(clock), .in1(R522));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op648 (.out1(R649), .clock(clock), .in1(R648));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op766 (.out1(R767), .clock(clock), .in1(R766));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op883 (.out1(R884), .clock(clock), .in1(R883));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op992 (.out1(R993), .clock(clock), .in1(R992));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1100 (.out1(R1101), .clock(clock), .in1(R1100));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1200 (.out1(R1201), .clock(clock), .in1(R1200));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1299 (.out1(R1300), .clock(clock), .in1(R1299));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1390 (.out1(R1391), .clock(clock), .in1(R1390));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1480 (.out1(R1481), .clock(clock), .in1(R1480));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1562 (.out1(R1563), .clock(clock), .in1(R1562));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1643 (.out1(R1644), .clock(clock), .in1(R1643));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1715 (.out1(R1716), .clock(clock), .in1(R1715));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1787 (.out1(R1788), .clock(clock), .in1(R1787));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1850 (.out1(R1851), .clock(clock), .in1(R1850));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1913 (.out1(R1914), .clock(clock), .in1(R1913));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1967 (.out1(R1968), .clock(clock), .in1(R1967));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2020 (.out1(R2021), .clock(clock), .in1(R2020));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2065 (.out1(R2066), .clock(clock), .in1(R2065));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2109 (.out1(R2110), .clock(clock), .in1(R2109));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2145 (.out1(R2146), .clock(clock), .in1(R2145));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2180 (.out1(R2181), .clock(clock), .in1(R2180));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2207 (.out1(R2208), .clock(clock), .in1(R2207));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2233 (.out1(R2234), .clock(clock), .in1(R2233));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2251 (.out1(R2252), .clock(clock), .in1(_160));
  SRAM op185 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_161),.ADR(R2252));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op396 (.out1(R397), .clock(clock), .in1(R396));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op523 (.out1(R524), .clock(clock), .in1(R523));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op649 (.out1(R650), .clock(clock), .in1(R649));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op767 (.out1(R768), .clock(clock), .in1(R767));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op884 (.out1(R885), .clock(clock), .in1(R884));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op993 (.out1(R994), .clock(clock), .in1(R993));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1101 (.out1(R1102), .clock(clock), .in1(R1101));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1201 (.out1(R1202), .clock(clock), .in1(R1201));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1300 (.out1(R1301), .clock(clock), .in1(R1300));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1391 (.out1(R1392), .clock(clock), .in1(R1391));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1481 (.out1(R1482), .clock(clock), .in1(R1481));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1563 (.out1(R1564), .clock(clock), .in1(R1563));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1644 (.out1(R1645), .clock(clock), .in1(R1644));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1716 (.out1(R1717), .clock(clock), .in1(R1716));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1788 (.out1(R1789), .clock(clock), .in1(R1788));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1851 (.out1(R1852), .clock(clock), .in1(R1851));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1914 (.out1(R1915), .clock(clock), .in1(R1914));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1968 (.out1(R1969), .clock(clock), .in1(R1968));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2021 (.out1(R2022), .clock(clock), .in1(R2021));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2066 (.out1(R2067), .clock(clock), .in1(R2066));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2110 (.out1(R2111), .clock(clock), .in1(R2110));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2146 (.out1(R2147), .clock(clock), .in1(R2146));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2181 (.out1(R2182), .clock(clock), .in1(R2181));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2208 (.out1(R2209), .clock(clock), .in1(R2208));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2234 (.out1(R2235), .clock(clock), .in1(R2234));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2252 (.out1(R2253), .clock(clock), .in1(_161));
  NE_EXPR #(.BITSIZE_in1(32), .BITSIZE_in2(1),.BITSIZE_out1(1)) op186 (.out1(ifout186), .in1(R2253), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op187 (.out1(_162), .in1(R2235));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op188 (.out1(_163), .in1(_162), .in2(2 'd 2));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op397 (.out1(R398), .clock(clock), .in1(R397));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op524 (.out1(R525), .clock(clock), .in1(R524));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op650 (.out1(R651), .clock(clock), .in1(R650));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op768 (.out1(R769), .clock(clock), .in1(R768));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op885 (.out1(R886), .clock(clock), .in1(R885));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op994 (.out1(R995), .clock(clock), .in1(R994));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1102 (.out1(R1103), .clock(clock), .in1(R1102));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1202 (.out1(R1203), .clock(clock), .in1(R1202));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1301 (.out1(R1302), .clock(clock), .in1(R1301));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1392 (.out1(R1393), .clock(clock), .in1(R1392));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1482 (.out1(R1483), .clock(clock), .in1(R1482));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1564 (.out1(R1565), .clock(clock), .in1(R1564));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1645 (.out1(R1646), .clock(clock), .in1(R1645));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1717 (.out1(R1718), .clock(clock), .in1(R1717));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1789 (.out1(R1790), .clock(clock), .in1(R1789));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1852 (.out1(R1853), .clock(clock), .in1(R1852));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1915 (.out1(R1916), .clock(clock), .in1(R1915));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1969 (.out1(R1970), .clock(clock), .in1(R1969));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2022 (.out1(R2023), .clock(clock), .in1(R2022));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2067 (.out1(R2068), .clock(clock), .in1(R2067));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2111 (.out1(R2112), .clock(clock), .in1(R2111));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2147 (.out1(R2148), .clock(clock), .in1(R2147));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2182 (.out1(R2183), .clock(clock), .in1(R2182));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2209 (.out1(R2210), .clock(clock), .in1(R2209));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2235 (.out1(R2236), .clock(clock), .in1(R2235));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2253 (.out1(R2254), .clock(clock), .in1(ifout186));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2270 (.out1(R2271), .clock(clock), .in1(_163));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op189 (.out1(_164), .in1(C112_281_D), .in2(R2271));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op398 (.out1(R399), .clock(clock), .in1(R398));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op525 (.out1(R526), .clock(clock), .in1(R525));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op651 (.out1(R652), .clock(clock), .in1(R651));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op769 (.out1(R770), .clock(clock), .in1(R769));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op886 (.out1(R887), .clock(clock), .in1(R886));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op995 (.out1(R996), .clock(clock), .in1(R995));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1103 (.out1(R1104), .clock(clock), .in1(R1103));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1203 (.out1(R1204), .clock(clock), .in1(R1203));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1302 (.out1(R1303), .clock(clock), .in1(R1302));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1393 (.out1(R1394), .clock(clock), .in1(R1393));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1483 (.out1(R1484), .clock(clock), .in1(R1483));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1565 (.out1(R1566), .clock(clock), .in1(R1565));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1646 (.out1(R1647), .clock(clock), .in1(R1646));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1718 (.out1(R1719), .clock(clock), .in1(R1718));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1790 (.out1(R1791), .clock(clock), .in1(R1790));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1853 (.out1(R1854), .clock(clock), .in1(R1853));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1916 (.out1(R1917), .clock(clock), .in1(R1916));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1970 (.out1(R1971), .clock(clock), .in1(R1970));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2023 (.out1(R2024), .clock(clock), .in1(R2023));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2068 (.out1(R2069), .clock(clock), .in1(R2068));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2112 (.out1(R2113), .clock(clock), .in1(R2112));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2148 (.out1(R2149), .clock(clock), .in1(R2148));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2183 (.out1(R2184), .clock(clock), .in1(R2183));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2210 (.out1(R2211), .clock(clock), .in1(R2210));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2236 (.out1(R2237), .clock(clock), .in1(R2236));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2254 (.out1(R2255), .clock(clock), .in1(R2254));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2271 (.out1(R2272), .clock(clock), .in1(_164));
  SRAM op190 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_165),.ADR(R2272));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op399 (.out1(R400), .clock(clock), .in1(R399));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op526 (.out1(R527), .clock(clock), .in1(R526));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op652 (.out1(R653), .clock(clock), .in1(R652));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op770 (.out1(R771), .clock(clock), .in1(R770));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op887 (.out1(R888), .clock(clock), .in1(R887));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op996 (.out1(R997), .clock(clock), .in1(R996));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1104 (.out1(R1105), .clock(clock), .in1(R1104));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1204 (.out1(R1205), .clock(clock), .in1(R1204));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1303 (.out1(R1304), .clock(clock), .in1(R1303));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1394 (.out1(R1395), .clock(clock), .in1(R1394));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1484 (.out1(R1485), .clock(clock), .in1(R1484));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1566 (.out1(R1567), .clock(clock), .in1(R1566));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1647 (.out1(R1648), .clock(clock), .in1(R1647));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1719 (.out1(R1720), .clock(clock), .in1(R1719));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1791 (.out1(R1792), .clock(clock), .in1(R1791));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1854 (.out1(R1855), .clock(clock), .in1(R1854));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1917 (.out1(R1918), .clock(clock), .in1(R1917));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1971 (.out1(R1972), .clock(clock), .in1(R1971));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2024 (.out1(R2025), .clock(clock), .in1(R2024));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2069 (.out1(R2070), .clock(clock), .in1(R2069));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2113 (.out1(R2114), .clock(clock), .in1(R2113));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2149 (.out1(R2150), .clock(clock), .in1(R2149));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2184 (.out1(R2185), .clock(clock), .in1(R2184));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2211 (.out1(R2212), .clock(clock), .in1(R2211));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2237 (.out1(R2238), .clock(clock), .in1(R2237));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2255 (.out1(R2256), .clock(clock), .in1(R2255));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2272 (.out1(R2273), .clock(clock), .in1(_165));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op191 (.out1(_166), .in1(R2273), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op400 (.out1(R401), .clock(clock), .in1(R400));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op527 (.out1(R528), .clock(clock), .in1(R527));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op653 (.out1(R654), .clock(clock), .in1(R653));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op771 (.out1(R772), .clock(clock), .in1(R771));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op888 (.out1(R889), .clock(clock), .in1(R888));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op997 (.out1(R998), .clock(clock), .in1(R997));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1105 (.out1(R1106), .clock(clock), .in1(R1105));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1205 (.out1(R1206), .clock(clock), .in1(R1205));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1304 (.out1(R1305), .clock(clock), .in1(R1304));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1395 (.out1(R1396), .clock(clock), .in1(R1395));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1485 (.out1(R1486), .clock(clock), .in1(R1485));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1567 (.out1(R1568), .clock(clock), .in1(R1567));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1648 (.out1(R1649), .clock(clock), .in1(R1648));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1720 (.out1(R1721), .clock(clock), .in1(R1720));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1792 (.out1(R1793), .clock(clock), .in1(R1792));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1855 (.out1(R1856), .clock(clock), .in1(R1855));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1918 (.out1(R1919), .clock(clock), .in1(R1918));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1972 (.out1(R1973), .clock(clock), .in1(R1972));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2025 (.out1(R2026), .clock(clock), .in1(R2025));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2070 (.out1(R2071), .clock(clock), .in1(R2070));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2114 (.out1(R2115), .clock(clock), .in1(R2114));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2150 (.out1(R2151), .clock(clock), .in1(R2150));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2185 (.out1(R2186), .clock(clock), .in1(R2185));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2212 (.out1(R2213), .clock(clock), .in1(R2212));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2238 (.out1(R2239), .clock(clock), .in1(R2238));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2256 (.out1(R2257), .clock(clock), .in1(R2256));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2273 (.out1(R2274), .clock(clock), .in1(_166));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(4), .BITSIZE_out1(32), .PRECISION(32)) op192 (.out1(_167), .in1(R2274), .in2(4 'd 8));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op401 (.out1(R402), .clock(clock), .in1(R401));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op528 (.out1(R529), .clock(clock), .in1(R528));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op654 (.out1(R655), .clock(clock), .in1(R654));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op772 (.out1(R773), .clock(clock), .in1(R772));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op889 (.out1(R890), .clock(clock), .in1(R889));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op998 (.out1(R999), .clock(clock), .in1(R998));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1106 (.out1(R1107), .clock(clock), .in1(R1106));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1206 (.out1(R1207), .clock(clock), .in1(R1206));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1305 (.out1(R1306), .clock(clock), .in1(R1305));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1396 (.out1(R1397), .clock(clock), .in1(R1396));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1486 (.out1(R1487), .clock(clock), .in1(R1486));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1568 (.out1(R1569), .clock(clock), .in1(R1568));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1649 (.out1(R1650), .clock(clock), .in1(R1649));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1721 (.out1(R1722), .clock(clock), .in1(R1721));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1793 (.out1(R1794), .clock(clock), .in1(R1793));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1856 (.out1(R1857), .clock(clock), .in1(R1856));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1919 (.out1(R1920), .clock(clock), .in1(R1919));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1973 (.out1(R1974), .clock(clock), .in1(R1973));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2026 (.out1(R2027), .clock(clock), .in1(R2026));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2071 (.out1(R2072), .clock(clock), .in1(R2071));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2115 (.out1(R2116), .clock(clock), .in1(R2115));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2151 (.out1(R2152), .clock(clock), .in1(R2151));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2186 (.out1(R2187), .clock(clock), .in1(R2186));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2213 (.out1(R2214), .clock(clock), .in1(R2213));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2239 (.out1(R2240), .clock(clock), .in1(R2239));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2257 (.out1(R2258), .clock(clock), .in1(R2257));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2274 (.out1(R2275), .clock(clock), .in1(_167));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(4), .BITSIZE_out1(64), .PRECISION(64)) op193 (.out1(_168), .in1(ip2_259_D), .in2(4 'd 8));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op194 (.out1(_169), .in1(_168));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(8), .BITSIZE_out1(32)) op195 (.out1(_170), .in1(_169), .in2(8 'd 255));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op196 (.out1(idx_284), .in1(R2275), .in2(_170));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op402 (.out1(R403), .clock(clock), .in1(R402));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op529 (.out1(R530), .clock(clock), .in1(R529));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op655 (.out1(R656), .clock(clock), .in1(R655));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op773 (.out1(R774), .clock(clock), .in1(R773));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op890 (.out1(R891), .clock(clock), .in1(R890));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op999 (.out1(R1000), .clock(clock), .in1(R999));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1107 (.out1(R1108), .clock(clock), .in1(R1107));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1207 (.out1(R1208), .clock(clock), .in1(R1207));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1306 (.out1(R1307), .clock(clock), .in1(R1306));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1397 (.out1(R1398), .clock(clock), .in1(R1397));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1487 (.out1(R1488), .clock(clock), .in1(R1487));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1569 (.out1(R1570), .clock(clock), .in1(R1569));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1650 (.out1(R1651), .clock(clock), .in1(R1650));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1722 (.out1(R1723), .clock(clock), .in1(R1722));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1794 (.out1(R1795), .clock(clock), .in1(R1794));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1857 (.out1(R1858), .clock(clock), .in1(R1857));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1920 (.out1(R1921), .clock(clock), .in1(R1920));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1974 (.out1(R1975), .clock(clock), .in1(R1974));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2027 (.out1(R2028), .clock(clock), .in1(R2027));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2072 (.out1(R2073), .clock(clock), .in1(R2072));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2116 (.out1(R2117), .clock(clock), .in1(R2116));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2152 (.out1(R2153), .clock(clock), .in1(R2152));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2187 (.out1(R2188), .clock(clock), .in1(R2187));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2214 (.out1(R2215), .clock(clock), .in1(R2214));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2240 (.out1(R2241), .clock(clock), .in1(R2240));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2258 (.out1(R2259), .clock(clock), .in1(R2258));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2275 (.out1(R2276), .clock(clock), .in1(idx_284));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op197 (.out1(_171), .in1(R2276));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op198 (.out1(_172), .in1(_171), .in2(2 'd 2));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op403 (.out1(R404), .clock(clock), .in1(R403));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op530 (.out1(R531), .clock(clock), .in1(R530));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op656 (.out1(R657), .clock(clock), .in1(R656));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op774 (.out1(R775), .clock(clock), .in1(R774));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op891 (.out1(R892), .clock(clock), .in1(R891));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1000 (.out1(R1001), .clock(clock), .in1(R1000));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1108 (.out1(R1109), .clock(clock), .in1(R1108));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1208 (.out1(R1209), .clock(clock), .in1(R1208));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1307 (.out1(R1308), .clock(clock), .in1(R1307));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1398 (.out1(R1399), .clock(clock), .in1(R1398));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1488 (.out1(R1489), .clock(clock), .in1(R1488));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1570 (.out1(R1571), .clock(clock), .in1(R1570));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1651 (.out1(R1652), .clock(clock), .in1(R1651));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1723 (.out1(R1724), .clock(clock), .in1(R1723));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1795 (.out1(R1796), .clock(clock), .in1(R1795));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1858 (.out1(R1859), .clock(clock), .in1(R1858));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1921 (.out1(R1922), .clock(clock), .in1(R1921));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1975 (.out1(R1976), .clock(clock), .in1(R1975));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2028 (.out1(R2029), .clock(clock), .in1(R2028));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2073 (.out1(R2074), .clock(clock), .in1(R2073));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2117 (.out1(R2118), .clock(clock), .in1(R2117));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2153 (.out1(R2154), .clock(clock), .in1(R2153));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2188 (.out1(R2189), .clock(clock), .in1(R2188));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2215 (.out1(R2216), .clock(clock), .in1(R2215));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2241 (.out1(R2242), .clock(clock), .in1(R2241));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2259 (.out1(R2260), .clock(clock), .in1(R2259));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2276 (.out1(R2277), .clock(clock), .in1(R2276));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2285 (.out1(R2286), .clock(clock), .in1(_172));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op199 (.out1(_173), .in1(C120_285_D), .in2(R2286));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op404 (.out1(R405), .clock(clock), .in1(R404));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op531 (.out1(R532), .clock(clock), .in1(R531));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op657 (.out1(R658), .clock(clock), .in1(R657));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op775 (.out1(R776), .clock(clock), .in1(R775));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op892 (.out1(R893), .clock(clock), .in1(R892));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1001 (.out1(R1002), .clock(clock), .in1(R1001));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1109 (.out1(R1110), .clock(clock), .in1(R1109));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1209 (.out1(R1210), .clock(clock), .in1(R1209));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1308 (.out1(R1309), .clock(clock), .in1(R1308));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1399 (.out1(R1400), .clock(clock), .in1(R1399));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1489 (.out1(R1490), .clock(clock), .in1(R1489));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1571 (.out1(R1572), .clock(clock), .in1(R1571));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1652 (.out1(R1653), .clock(clock), .in1(R1652));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1724 (.out1(R1725), .clock(clock), .in1(R1724));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1796 (.out1(R1797), .clock(clock), .in1(R1796));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1859 (.out1(R1860), .clock(clock), .in1(R1859));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1922 (.out1(R1923), .clock(clock), .in1(R1922));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1976 (.out1(R1977), .clock(clock), .in1(R1976));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2029 (.out1(R2030), .clock(clock), .in1(R2029));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2074 (.out1(R2075), .clock(clock), .in1(R2074));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2118 (.out1(R2119), .clock(clock), .in1(R2118));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2154 (.out1(R2155), .clock(clock), .in1(R2154));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2189 (.out1(R2190), .clock(clock), .in1(R2189));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2216 (.out1(R2217), .clock(clock), .in1(R2216));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2242 (.out1(R2243), .clock(clock), .in1(R2242));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2260 (.out1(R2261), .clock(clock), .in1(R2260));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2277 (.out1(R2278), .clock(clock), .in1(R2277));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2286 (.out1(R2287), .clock(clock), .in1(_173));
  SRAM op200 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_174),.ADR(R2287));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op405 (.out1(R406), .clock(clock), .in1(R405));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op532 (.out1(R533), .clock(clock), .in1(R532));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op658 (.out1(R659), .clock(clock), .in1(R658));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op776 (.out1(R777), .clock(clock), .in1(R776));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op893 (.out1(R894), .clock(clock), .in1(R893));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1002 (.out1(R1003), .clock(clock), .in1(R1002));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1110 (.out1(R1111), .clock(clock), .in1(R1110));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1210 (.out1(R1211), .clock(clock), .in1(R1210));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1309 (.out1(R1310), .clock(clock), .in1(R1309));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1400 (.out1(R1401), .clock(clock), .in1(R1400));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1490 (.out1(R1491), .clock(clock), .in1(R1490));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1572 (.out1(R1573), .clock(clock), .in1(R1572));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1653 (.out1(R1654), .clock(clock), .in1(R1653));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1725 (.out1(R1726), .clock(clock), .in1(R1725));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1797 (.out1(R1798), .clock(clock), .in1(R1797));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1860 (.out1(R1861), .clock(clock), .in1(R1860));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1923 (.out1(R1924), .clock(clock), .in1(R1923));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1977 (.out1(R1978), .clock(clock), .in1(R1977));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2030 (.out1(R2031), .clock(clock), .in1(R2030));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2075 (.out1(R2076), .clock(clock), .in1(R2075));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2119 (.out1(R2120), .clock(clock), .in1(R2119));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2155 (.out1(R2156), .clock(clock), .in1(R2155));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2190 (.out1(R2191), .clock(clock), .in1(R2190));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2217 (.out1(R2218), .clock(clock), .in1(R2217));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2243 (.out1(R2244), .clock(clock), .in1(R2243));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2261 (.out1(R2262), .clock(clock), .in1(R2261));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2278 (.out1(R2279), .clock(clock), .in1(R2278));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2287 (.out1(R2288), .clock(clock), .in1(_174));
  NE_EXPR #(.BITSIZE_in1(32), .BITSIZE_in2(1),.BITSIZE_out1(1)) op201 (.out1(ifout201), .in1(R2288), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op202 (.out1(_175), .in1(R2279));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op203 (.out1(_176), .in1(_175), .in2(2 'd 2));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op406 (.out1(R407), .clock(clock), .in1(R406));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op533 (.out1(R534), .clock(clock), .in1(R533));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op659 (.out1(R660), .clock(clock), .in1(R659));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op777 (.out1(R778), .clock(clock), .in1(R777));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op894 (.out1(R895), .clock(clock), .in1(R894));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1003 (.out1(R1004), .clock(clock), .in1(R1003));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1111 (.out1(R1112), .clock(clock), .in1(R1111));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1211 (.out1(R1212), .clock(clock), .in1(R1211));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1310 (.out1(R1311), .clock(clock), .in1(R1310));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1401 (.out1(R1402), .clock(clock), .in1(R1401));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1491 (.out1(R1492), .clock(clock), .in1(R1491));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1573 (.out1(R1574), .clock(clock), .in1(R1573));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1654 (.out1(R1655), .clock(clock), .in1(R1654));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1726 (.out1(R1727), .clock(clock), .in1(R1726));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1798 (.out1(R1799), .clock(clock), .in1(R1798));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1861 (.out1(R1862), .clock(clock), .in1(R1861));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1924 (.out1(R1925), .clock(clock), .in1(R1924));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1978 (.out1(R1979), .clock(clock), .in1(R1978));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2031 (.out1(R2032), .clock(clock), .in1(R2031));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2076 (.out1(R2077), .clock(clock), .in1(R2076));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2120 (.out1(R2121), .clock(clock), .in1(R2120));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2156 (.out1(R2157), .clock(clock), .in1(R2156));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2191 (.out1(R2192), .clock(clock), .in1(R2191));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2218 (.out1(R2219), .clock(clock), .in1(R2218));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2244 (.out1(R2245), .clock(clock), .in1(R2244));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2262 (.out1(R2263), .clock(clock), .in1(R2262));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2279 (.out1(R2280), .clock(clock), .in1(R2279));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2288 (.out1(R2289), .clock(clock), .in1(ifout201));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2296 (.out1(R2297), .clock(clock), .in1(_176));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op204 (.out1(_177), .in1(C120_285_D), .in2(R2297));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op407 (.out1(R408), .clock(clock), .in1(R407));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op534 (.out1(R535), .clock(clock), .in1(R534));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op660 (.out1(R661), .clock(clock), .in1(R660));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op778 (.out1(R779), .clock(clock), .in1(R778));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op895 (.out1(R896), .clock(clock), .in1(R895));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1004 (.out1(R1005), .clock(clock), .in1(R1004));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1112 (.out1(R1113), .clock(clock), .in1(R1112));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1212 (.out1(R1213), .clock(clock), .in1(R1212));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1311 (.out1(R1312), .clock(clock), .in1(R1311));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1402 (.out1(R1403), .clock(clock), .in1(R1402));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1492 (.out1(R1493), .clock(clock), .in1(R1492));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1574 (.out1(R1575), .clock(clock), .in1(R1574));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1655 (.out1(R1656), .clock(clock), .in1(R1655));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1727 (.out1(R1728), .clock(clock), .in1(R1727));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1799 (.out1(R1800), .clock(clock), .in1(R1799));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1862 (.out1(R1863), .clock(clock), .in1(R1862));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1925 (.out1(R1926), .clock(clock), .in1(R1925));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1979 (.out1(R1980), .clock(clock), .in1(R1979));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2032 (.out1(R2033), .clock(clock), .in1(R2032));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2077 (.out1(R2078), .clock(clock), .in1(R2077));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2121 (.out1(R2122), .clock(clock), .in1(R2121));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2157 (.out1(R2158), .clock(clock), .in1(R2157));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2192 (.out1(R2193), .clock(clock), .in1(R2192));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2219 (.out1(R2220), .clock(clock), .in1(R2219));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2245 (.out1(R2246), .clock(clock), .in1(R2245));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2263 (.out1(R2264), .clock(clock), .in1(R2263));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2280 (.out1(R2281), .clock(clock), .in1(R2280));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2289 (.out1(R2290), .clock(clock), .in1(R2289));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2297 (.out1(R2298), .clock(clock), .in1(_177));
  SRAM op205 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_178),.ADR(R2298));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op408 (.out1(R409), .clock(clock), .in1(R408));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op535 (.out1(R536), .clock(clock), .in1(R535));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op661 (.out1(R662), .clock(clock), .in1(R661));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op779 (.out1(R780), .clock(clock), .in1(R779));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op896 (.out1(R897), .clock(clock), .in1(R896));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1005 (.out1(R1006), .clock(clock), .in1(R1005));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1113 (.out1(R1114), .clock(clock), .in1(R1113));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1213 (.out1(R1214), .clock(clock), .in1(R1213));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1312 (.out1(R1313), .clock(clock), .in1(R1312));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1403 (.out1(R1404), .clock(clock), .in1(R1403));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1493 (.out1(R1494), .clock(clock), .in1(R1493));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1575 (.out1(R1576), .clock(clock), .in1(R1575));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1656 (.out1(R1657), .clock(clock), .in1(R1656));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1728 (.out1(R1729), .clock(clock), .in1(R1728));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1800 (.out1(R1801), .clock(clock), .in1(R1800));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1863 (.out1(R1864), .clock(clock), .in1(R1863));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1926 (.out1(R1927), .clock(clock), .in1(R1926));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1980 (.out1(R1981), .clock(clock), .in1(R1980));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2033 (.out1(R2034), .clock(clock), .in1(R2033));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2078 (.out1(R2079), .clock(clock), .in1(R2078));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2122 (.out1(R2123), .clock(clock), .in1(R2122));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2158 (.out1(R2159), .clock(clock), .in1(R2158));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2193 (.out1(R2194), .clock(clock), .in1(R2193));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2220 (.out1(R2221), .clock(clock), .in1(R2220));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2246 (.out1(R2247), .clock(clock), .in1(R2246));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2264 (.out1(R2265), .clock(clock), .in1(R2264));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2281 (.out1(R2282), .clock(clock), .in1(R2281));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2290 (.out1(R2291), .clock(clock), .in1(R2290));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2298 (.out1(R2299), .clock(clock), .in1(_178));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op206 (.out1(_179), .in1(R2299), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op409 (.out1(R410), .clock(clock), .in1(R409));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op536 (.out1(R537), .clock(clock), .in1(R536));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op662 (.out1(R663), .clock(clock), .in1(R662));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op780 (.out1(R781), .clock(clock), .in1(R780));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op897 (.out1(R898), .clock(clock), .in1(R897));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1006 (.out1(R1007), .clock(clock), .in1(R1006));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1114 (.out1(R1115), .clock(clock), .in1(R1114));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1214 (.out1(R1215), .clock(clock), .in1(R1214));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1313 (.out1(R1314), .clock(clock), .in1(R1313));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1404 (.out1(R1405), .clock(clock), .in1(R1404));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1494 (.out1(R1495), .clock(clock), .in1(R1494));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1576 (.out1(R1577), .clock(clock), .in1(R1576));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1657 (.out1(R1658), .clock(clock), .in1(R1657));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1729 (.out1(R1730), .clock(clock), .in1(R1729));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1801 (.out1(R1802), .clock(clock), .in1(R1801));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1864 (.out1(R1865), .clock(clock), .in1(R1864));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1927 (.out1(R1928), .clock(clock), .in1(R1927));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1981 (.out1(R1982), .clock(clock), .in1(R1981));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2034 (.out1(R2035), .clock(clock), .in1(R2034));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2079 (.out1(R2080), .clock(clock), .in1(R2079));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2123 (.out1(R2124), .clock(clock), .in1(R2123));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2159 (.out1(R2160), .clock(clock), .in1(R2159));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2194 (.out1(R2195), .clock(clock), .in1(R2194));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2221 (.out1(R2222), .clock(clock), .in1(R2221));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2247 (.out1(R2248), .clock(clock), .in1(R2247));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2265 (.out1(R2266), .clock(clock), .in1(R2265));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2282 (.out1(R2283), .clock(clock), .in1(R2282));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2291 (.out1(R2292), .clock(clock), .in1(R2291));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2299 (.out1(R2300), .clock(clock), .in1(_179));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(4), .BITSIZE_out1(32), .PRECISION(32)) op207 (.out1(_180), .in1(R2300), .in2(4 'd 8));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op410 (.out1(R411), .clock(clock), .in1(R410));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op537 (.out1(R538), .clock(clock), .in1(R537));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op663 (.out1(R664), .clock(clock), .in1(R663));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op781 (.out1(R782), .clock(clock), .in1(R781));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op898 (.out1(R899), .clock(clock), .in1(R898));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1007 (.out1(R1008), .clock(clock), .in1(R1007));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1115 (.out1(R1116), .clock(clock), .in1(R1115));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1215 (.out1(R1216), .clock(clock), .in1(R1215));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1314 (.out1(R1315), .clock(clock), .in1(R1314));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1405 (.out1(R1406), .clock(clock), .in1(R1405));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1495 (.out1(R1496), .clock(clock), .in1(R1495));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1577 (.out1(R1578), .clock(clock), .in1(R1577));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1658 (.out1(R1659), .clock(clock), .in1(R1658));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1730 (.out1(R1731), .clock(clock), .in1(R1730));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1802 (.out1(R1803), .clock(clock), .in1(R1802));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1865 (.out1(R1866), .clock(clock), .in1(R1865));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1928 (.out1(R1929), .clock(clock), .in1(R1928));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1982 (.out1(R1983), .clock(clock), .in1(R1982));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2035 (.out1(R2036), .clock(clock), .in1(R2035));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2080 (.out1(R2081), .clock(clock), .in1(R2080));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2124 (.out1(R2125), .clock(clock), .in1(R2124));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2160 (.out1(R2161), .clock(clock), .in1(R2160));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2195 (.out1(R2196), .clock(clock), .in1(R2195));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2222 (.out1(R2223), .clock(clock), .in1(R2222));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2248 (.out1(R2249), .clock(clock), .in1(R2248));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2266 (.out1(R2267), .clock(clock), .in1(R2266));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2283 (.out1(R2284), .clock(clock), .in1(R2283));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2292 (.out1(R2293), .clock(clock), .in1(R2292));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2300 (.out1(R2301), .clock(clock), .in1(_180));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op208 (.out1(_181), .in1(ip2_259_D));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(8), .BITSIZE_out1(32)) op209 (.out1(_182), .in1(_181), .in2(8 'd 255));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op210 (.out1(idx_288), .in1(R2301), .in2(_182));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op411 (.out1(R412), .clock(clock), .in1(R411));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op538 (.out1(R539), .clock(clock), .in1(R538));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op664 (.out1(R665), .clock(clock), .in1(R664));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op782 (.out1(R783), .clock(clock), .in1(R782));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op899 (.out1(R900), .clock(clock), .in1(R899));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1008 (.out1(R1009), .clock(clock), .in1(R1008));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1116 (.out1(R1117), .clock(clock), .in1(R1116));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1216 (.out1(R1217), .clock(clock), .in1(R1216));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1315 (.out1(R1316), .clock(clock), .in1(R1315));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1406 (.out1(R1407), .clock(clock), .in1(R1406));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1496 (.out1(R1497), .clock(clock), .in1(R1496));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1578 (.out1(R1579), .clock(clock), .in1(R1578));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1659 (.out1(R1660), .clock(clock), .in1(R1659));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1731 (.out1(R1732), .clock(clock), .in1(R1731));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1803 (.out1(R1804), .clock(clock), .in1(R1803));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1866 (.out1(R1867), .clock(clock), .in1(R1866));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1929 (.out1(R1930), .clock(clock), .in1(R1929));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1983 (.out1(R1984), .clock(clock), .in1(R1983));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2036 (.out1(R2037), .clock(clock), .in1(R2036));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2081 (.out1(R2082), .clock(clock), .in1(R2081));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2125 (.out1(R2126), .clock(clock), .in1(R2125));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2161 (.out1(R2162), .clock(clock), .in1(R2161));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2196 (.out1(R2197), .clock(clock), .in1(R2196));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2223 (.out1(R2224), .clock(clock), .in1(R2223));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2249 (.out1(R2250), .clock(clock), .in1(R2249));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2267 (.out1(R2268), .clock(clock), .in1(R2267));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2284 (.out1(R2285), .clock(clock), .in1(R2284));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2293 (.out1(R2294), .clock(clock), .in1(R2293));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2301 (.out1(R2302), .clock(clock), .in1(idx_288));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op243 (.out1(_207), .in1(R1660));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op239 (.out1(_204), .in1(R1804));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op235 (.out1(_201), .in1(R1930));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op231 (.out1(_198), .in1(R2037));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op227 (.out1(_195), .in1(R2126));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op223 (.out1(_192), .in1(R2197));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op219 (.out1(_189), .in1(R2250));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op215 (.out1(_186), .in1(R2285));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op211 (.out1(_183), .in1(R2302));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op244 (.out1(_208), .in1(N64_257_D), .in2(_207));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op240 (.out1(_205), .in1(N72_262_D), .in2(_204));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op236 (.out1(_202), .in1(N80_266_D), .in2(_201));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op232 (.out1(_199), .in1(N88_270_D), .in2(_198));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op228 (.out1(_196), .in1(N96_274_D), .in2(_195));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op224 (.out1(_193), .in1(N104_278_D), .in2(_192));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op220 (.out1(_190), .in1(N112_282_D), .in2(_189));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op216 (.out1(_187), .in1(N120_286_D), .in2(_186));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op212 (.out1(_184), .in1(N128_289_D), .in2(_183));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op412 (.out1(R413), .clock(clock), .in1(R412));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op539 (.out1(R540), .clock(clock), .in1(R539));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op665 (.out1(R666), .clock(clock), .in1(R665));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op783 (.out1(R784), .clock(clock), .in1(R783));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op900 (.out1(R901), .clock(clock), .in1(R900));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1009 (.out1(R1010), .clock(clock), .in1(R1009));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1117 (.out1(R1118), .clock(clock), .in1(R1117));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1217 (.out1(R1218), .clock(clock), .in1(R1217));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1316 (.out1(R1317), .clock(clock), .in1(R1316));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1407 (.out1(R1408), .clock(clock), .in1(R1407));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op1497 (.out1(R1498), .clock(clock), .in1(R1497));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1579 (.out1(R1580), .clock(clock), .in1(R1579));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1732 (.out1(R1733), .clock(clock), .in1(R1732));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1867 (.out1(R1868), .clock(clock), .in1(R1867));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1984 (.out1(R1985), .clock(clock), .in1(R1984));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2082 (.out1(R2083), .clock(clock), .in1(R2082));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2162 (.out1(R2163), .clock(clock), .in1(R2162));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2224 (.out1(R2225), .clock(clock), .in1(R2224));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2268 (.out1(R2269), .clock(clock), .in1(R2268));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2294 (.out1(R2295), .clock(clock), .in1(R2294));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2302 (.out1(R2303), .clock(clock), .in1(_208));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2303 (.out1(R2304), .clock(clock), .in1(_205));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2304 (.out1(R2305), .clock(clock), .in1(_202));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2305 (.out1(R2306), .clock(clock), .in1(_199));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2306 (.out1(R2307), .clock(clock), .in1(_196));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2307 (.out1(R2308), .clock(clock), .in1(_193));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2308 (.out1(R2309), .clock(clock), .in1(_190));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2309 (.out1(R2310), .clock(clock), .in1(_187));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2310 (.out1(R2311), .clock(clock), .in1(_184));
  SRAM op245 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_209),.ADR(R2303));
  SRAM op241 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_206),.ADR(R2304));
  SRAM op237 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_203),.ADR(R2305));
  SRAM op233 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_200),.ADR(R2306));
  SRAM op229 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_197),.ADR(R2307));
  SRAM op225 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_194),.ADR(R2308));
  SRAM op221 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_191),.ADR(R2309));
  SRAM op217 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_188),.ADR(R2310));
  SRAM op213 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_185),.ADR(R2311));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op267 (.out1(_225), .in1(R413));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op263 (.out1(_222), .in1(R666));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op259 (.out1(_219), .in1(R901));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op255 (.out1(_216), .in1(R1118));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op251 (.out1(_213), .in1(R1317));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op247 (.out1(_210), .in1(R1498));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op268 (.out1(_226), .in1(N16_233_D), .in2(_225));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op264 (.out1(_223), .in1(N24_237_D), .in2(_222));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op260 (.out1(_220), .in1(N32_241_D), .in2(_219));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op256 (.out1(_217), .in1(N40_245_D), .in2(_216));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op252 (.out1(_214), .in1(N48_249_D), .in2(_213));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op248 (.out1(_211), .in1(N56_253_D), .in2(_210));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op540 (.out1(R541), .clock(clock), .in1(R540));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op784 (.out1(R785), .clock(clock), .in1(R784));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1010 (.out1(R1011), .clock(clock), .in1(R1010));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1218 (.out1(R1219), .clock(clock), .in1(R1218));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1408 (.out1(R1409), .clock(clock), .in1(R1408));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1580 (.out1(R1581), .clock(clock), .in1(R1580));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1733 (.out1(R1734), .clock(clock), .in1(R1733));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1868 (.out1(R1869), .clock(clock), .in1(R1868));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1985 (.out1(R1986), .clock(clock), .in1(R1985));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2083 (.out1(R2084), .clock(clock), .in1(R2083));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2163 (.out1(R2164), .clock(clock), .in1(R2163));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2225 (.out1(R2226), .clock(clock), .in1(R2225));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2269 (.out1(R2270), .clock(clock), .in1(R2269));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op2295 (.out1(R2296), .clock(clock), .in1(R2295));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op2311 (.out1(R2312), .clock(clock), .in1(_209));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op2312 (.out1(R2313), .clock(clock), .in1(_206));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op2313 (.out1(R2314), .clock(clock), .in1(_203));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op2314 (.out1(R2315), .clock(clock), .in1(_200));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op2315 (.out1(R2316), .clock(clock), .in1(_197));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op2316 (.out1(R2317), .clock(clock), .in1(_194));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op2317 (.out1(R2318), .clock(clock), .in1(_191));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op2318 (.out1(R2319), .clock(clock), .in1(_188));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op2319 (.out1(R2320), .clock(clock), .in1(_185));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2320 (.out1(R2321), .clock(clock), .in1(_226));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2321 (.out1(R2322), .clock(clock), .in1(_223));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2322 (.out1(R2323), .clock(clock), .in1(_220));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2323 (.out1(R2324), .clock(clock), .in1(_217));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2324 (.out1(R2325), .clock(clock), .in1(_214));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2325 (.out1(R2326), .clock(clock), .in1(_211));
  SRAM op269 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_227),.ADR(R2321));
  SRAM op265 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_224),.ADR(R2322));
  SRAM op261 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_221),.ADR(R2323));
  SRAM op257 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_218),.ADR(R2324));
  SRAM op253 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_215),.ADR(R2325));
  SRAM op249 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_212),.ADR(R2326));
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op218 (.out1(_287), .in1(R2319));
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op214 (.out1(_290), .in1(R2320));
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op222 (.out1(_283), .in1(R2318));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op271 (.out1(mux0), .in1(_287), .in2(_290), .sel(R2296));
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op226 (.out1(_279), .in1(R2317));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op272 (.out1(mux1), .in1(_283), .in2(mux0), .sel(R2270));
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op230 (.out1(_275), .in1(R2316));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op273 (.out1(mux2), .in1(_279), .in2(mux1), .sel(R2226));
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op234 (.out1(_271), .in1(R2315));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op274 (.out1(mux3), .in1(_275), .in2(mux2), .sel(R2164));
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op238 (.out1(_267), .in1(R2314));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op275 (.out1(mux4), .in1(_271), .in2(mux3), .sel(R2084));
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op246 (.out1(_258), .in1(R2312));
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op242 (.out1(_263), .in1(R2313));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op276 (.out1(mux5), .in1(_267), .in2(mux4), .sel(R1986));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op541 (.out1(R542), .clock(clock), .in1(R541));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op785 (.out1(R786), .clock(clock), .in1(R785));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1011 (.out1(R1012), .clock(clock), .in1(R1011));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1219 (.out1(R1220), .clock(clock), .in1(R1219));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1409 (.out1(R1410), .clock(clock), .in1(R1409));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1581 (.out1(R1582), .clock(clock), .in1(R1581));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1734 (.out1(R1735), .clock(clock), .in1(R1734));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op1869 (.out1(R1870), .clock(clock), .in1(R1869));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op2326 (.out1(R2327), .clock(clock), .in1(_227));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op2327 (.out1(R2328), .clock(clock), .in1(_224));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op2328 (.out1(R2329), .clock(clock), .in1(_221));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op2329 (.out1(R2330), .clock(clock), .in1(_218));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op2330 (.out1(R2331), .clock(clock), .in1(_215));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op2331 (.out1(R2332), .clock(clock), .in1(_212));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op2332 (.out1(R2333), .clock(clock), .in1(_258));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op2333 (.out1(R2334), .clock(clock), .in1(_263));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op2334 (.out1(R2335), .clock(clock), .in1(mux5));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op277 (.out1(mux6), .in1(R2334), .in2(R2335), .sel(R1870));
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op250 (.out1(_254), .in1(R2332));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op278 (.out1(mux7), .in1(R2333), .in2(mux6), .sel(R1735));
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op254 (.out1(_250), .in1(R2331));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op279 (.out1(mux8), .in1(_254), .in2(mux7), .sel(R1582));
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op258 (.out1(_246), .in1(R2330));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op280 (.out1(mux9), .in1(_250), .in2(mux8), .sel(R1410));
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op262 (.out1(_242), .in1(R2329));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op281 (.out1(mux10), .in1(_246), .in2(mux9), .sel(R1220));
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op266 (.out1(_238), .in1(R2328));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op282 (.out1(mux11), .in1(_242), .in2(mux10), .sel(R1012));
  cast #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op270 (.out1(_234), .in1(R2327));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op283 (.out1(mux12), .in1(_238), .in2(mux11), .sel(R786));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op284 (.out1(mux13), .in1(_234), .in2(mux12), .sel(R542));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op2335 (.out1(R2336), .clock(clock), .in1(mux13));
endmodule