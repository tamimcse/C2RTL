`include "module_library.v"
`include "macros.v"

`timescale 1ns / 1ps
module top(clock, b16_popcnt_2529_D, b16_bitmap_2528_D, b24_popcnt_2540_D, b24_bitmap_2539_D, b32_popcnt_2550_D, b32_bitmap_2549_D, b40_popcnt_2560_D, b40_bitmap_2559_D, b48_popcnt_2570_D, b48_bitmap_2569_D, b56_popcnt_2580_D, b56_bitmap_2579_D, b64_popcnt_2590_D, b64_bitmap_2589_D, b72_popcnt_2601_D, b72_bitmap_2600_D, b80_popcnt_2611_D, b80_bitmap_2610_D, b88_popcnt_2621_D, b88_bitmap_2620_D, b96_popcnt_2631_D, b96_bitmap_2630_D, b104_popcnt_2641_D, b104_bitmap_2640_D, b112_popcnt_2651_D, b112_bitmap_2650_D, b120_popcnt_2661_D, b120_bitmap_2660_D, leafN_2531_D, b128_popcnt_2670_D, b128_bitmap_2669_D, c120_popcnt_2664_D, c120_bitmap_2659_D, c112_popcnt_2654_D, c112_bitmap_2649_D, c104_popcnt_2644_D, c104_bitmap_2639_D, c96_popcnt_2634_D, c96_bitmap_2629_D, c88_popcnt_2624_D, c88_bitmap_2619_D, c80_popcnt_2614_D, c80_bitmap_2609_D, c72_popcnt_2604_D, c72_bitmap_2599_D, ip2_2595_D, c64_popcnt_2593_D, c64_bitmap_2588_D, c56_popcnt_2583_D, c56_bitmap_2578_D, c48_popcnt_2573_D, c48_bitmap_2568_D, c40_popcnt_2563_D, c40_bitmap_2558_D, c32_popcnt_2553_D, c32_bitmap_2548_D, c24_popcnt_2543_D, c24_bitmap_2538_D, c16_popcnt_2533_D, c16_bitmap_2526_D, ip1_2522_D, R9124);
  //IN
  input clock;
  input [63:0] b16_popcnt_2529_D;
  input [63:0] b16_bitmap_2528_D;
  input [63:0] b24_popcnt_2540_D;
  input [63:0] b24_bitmap_2539_D;
  input [63:0] b32_popcnt_2550_D;
  input [63:0] b32_bitmap_2549_D;
  input [63:0] b40_popcnt_2560_D;
  input [63:0] b40_bitmap_2559_D;
  input [63:0] b48_popcnt_2570_D;
  input [63:0] b48_bitmap_2569_D;
  input [63:0] b56_popcnt_2580_D;
  input [63:0] b56_bitmap_2579_D;
  input [63:0] b64_popcnt_2590_D;
  input [63:0] b64_bitmap_2589_D;
  input [63:0] b72_popcnt_2601_D;
  input [63:0] b72_bitmap_2600_D;
  input [63:0] b80_popcnt_2611_D;
  input [63:0] b80_bitmap_2610_D;
  input [63:0] b88_popcnt_2621_D;
  input [63:0] b88_bitmap_2620_D;
  input [63:0] b96_popcnt_2631_D;
  input [63:0] b96_bitmap_2630_D;
  input [63:0] b104_popcnt_2641_D;
  input [63:0] b104_bitmap_2640_D;
  input [63:0] b112_popcnt_2651_D;
  input [63:0] b112_bitmap_2650_D;
  input [63:0] b120_popcnt_2661_D;
  input [63:0] b120_bitmap_2660_D;
  input [63:0] leafN_2531_D;
  input [63:0] b128_popcnt_2670_D;
  input [63:0] b128_bitmap_2669_D;
  input [63:0] c120_popcnt_2664_D;
  input [63:0] c120_bitmap_2659_D;
  input [63:0] c112_popcnt_2654_D;
  input [63:0] c112_bitmap_2649_D;
  input [63:0] c104_popcnt_2644_D;
  input [63:0] c104_bitmap_2639_D;
  input [63:0] c96_popcnt_2634_D;
  input [63:0] c96_bitmap_2629_D;
  input [63:0] c88_popcnt_2624_D;
  input [63:0] c88_bitmap_2619_D;
  input [63:0] c80_popcnt_2614_D;
  input [63:0] c80_bitmap_2609_D;
  input [63:0] c72_popcnt_2604_D;
  input [63:0] c72_bitmap_2599_D;
  input [63:0] ip2_2595_D;
  input [63:0] c64_popcnt_2593_D;
  input [63:0] c64_bitmap_2588_D;
  input [63:0] c56_popcnt_2583_D;
  input [63:0] c56_bitmap_2578_D;
  input [63:0] c48_popcnt_2573_D;
  input [63:0] c48_bitmap_2568_D;
  input [63:0] c40_popcnt_2563_D;
  input [63:0] c40_bitmap_2558_D;
  input [63:0] c32_popcnt_2553_D;
  input [63:0] c32_bitmap_2548_D;
  input [63:0] c24_popcnt_2543_D;
  input [63:0] c24_bitmap_2538_D;
  input [63:0] c16_popcnt_2533_D;
  input [63:0] c16_bitmap_2526_D;
  input [63:0] ip1_2522_D;
  //OUT
  output [7:0] R9124;
  //WIRES
  wire [7:0] R9124;
  wire [7:0] R9123;
  wire [7:0] R9122;
  wire [7:0] R9121;
  wire [7:0] R9120;
  wire [7:0] R9119;
  wire [7:0] R9118;
  wire [7:0] R9117;
  wire [7:0] R9116;
  wire [7:0] R9115;
  wire [7:0] R9114;
  wire [63:0] R9113;
  wire [63:0] R9112;
  wire [63:0] R9111;
  wire [63:0] R9110;
  wire [63:0] R9109;
  wire [63:0] R9108;
  wire [7:0] R9107;
  wire [7:0] R9106;
  wire [7:0] R9105;
  wire [7:0] R9104;
  wire [7:0] R9103;
  wire [7:0] R9102;
  wire [7:0] R9101;
  wire [7:0] R9100;
  wire [7:0] R9099;
  wire [31:0] R9098;
  wire [31:0] R9097;
  wire [31:0] R9096;
  wire [31:0] R9095;
  wire [31:0] R9094;
  wire [31:0] R9093;
  wire [63:0] R9092;
  wire [63:0] R9091;
  wire [63:0] R9090;
  wire [63:0] R9089;
  wire [63:0] R9088;
  wire [63:0] R9087;
  wire [63:0] R9086;
  wire [63:0] R9085;
  wire [63:0] R9084;
  wire [31:0] R9083;
  wire [31:0] R9082;
  wire [31:0] R9081;
  wire [31:0] R9080;
  wire [31:0] R9079;
  wire [31:0] R9078;
  wire [31:0] R9077;
  wire [31:0] R9076;
  wire [31:0] R9075;
  wire [63:0] R9074;
  wire [63:0] R9073;
  wire [63:0] R9072;
  wire [63:0] R9071;
  wire [63:0] R9070;
  wire [63:0] R9069;
  wire [31:0] R9068;
  wire [31:0] R9067;
  wire [31:0] R9066;
  wire [31:0] R9065;
  wire [31:0] R9064;
  wire [31:0] R9063;
  wire [63:0] R9062;
  wire [63:0] R9061;
  wire [63:0] R9060;
  wire [63:0] R9059;
  wire [63:0] R9058;
  wire [63:0] R9057;
  wire [63:0] R9056;
  wire [63:0] R9055;
  wire [63:0] R9054;
  wire [63:0] R9053;
  wire [63:0] R9052;
  wire [63:0] R9051;
  wire [63:0] R9050;
  wire [63:0] R9049;
  wire [63:0] R9048;
  wire [63:0] R9047;
  wire [63:0] R9046;
  wire [63:0] R9045;
  wire [63:0] R9044;
  wire [63:0] R9043;
  wire [63:0] R9042;
  wire [31:0] R9041;
  wire [31:0] R9040;
  wire [31:0] R9039;
  wire [31:0] R9038;
  wire [31:0] R9037;
  wire [31:0] R9036;
  wire [31:0] R9035;
  wire [31:0] R9034;
  wire [31:0] R9033;
  wire [63:0] R9032;
  wire [63:0] R9031;
  wire [63:0] R9030;
  wire [63:0] R9029;
  wire [63:0] R9028;
  wire [63:0] R9027;
  wire [63:0] R9026;
  wire [63:0] R9025;
  wire [63:0] R9024;
  wire [63:0] R9023;
  wire [63:0] R9022;
  wire [63:0] R9021;
  wire [63:0] R9020;
  wire [63:0] R9019;
  wire [63:0] R9018;
  wire [63:0] R9017;
  wire [63:0] R9016;
  wire [63:0] R9015;
  wire [63:0] R9014;
  wire [63:0] R9013;
  wire [63:0] R9012;
  wire [63:0] R9011;
  wire [63:0] R9010;
  wire [63:0] R9009;
  wire [63:0] R9008;
  wire [63:0] R9007;
  wire [63:0] R9006;
  wire [63:0] R9005;
  wire [63:0] R9004;
  wire [63:0] R9003;
  wire [63:0] R9002;
  wire [63:0] R9001;
  wire [63:0] R9000;
  wire [63:0] R8999;
  wire [63:0] R8998;
  wire [63:0] R8997;
  wire [63:0] R8996;
  wire [63:0] R8995;
  wire [63:0] R8994;
  wire [63:0] R8993;
  wire [63:0] R8992;
  wire [63:0] R8991;
  wire [63:0] R8990;
  wire [63:0] R8989;
  wire [63:0] R8988;
  wire [63:0] R8987;
  wire [63:0] R8986;
  wire [63:0] R8985;
  wire [63:0] R8984;
  wire [63:0] R8983;
  wire [63:0] R8982;
  wire [63:0] R8981;
  wire [63:0] R8980;
  wire [63:0] R8979;
  wire [63:0] R8978;
  wire [63:0] R8977;
  wire [63:0] R8976;
  wire [63:0] R8975;
  wire [63:0] R8974;
  wire [63:0] R8973;
  wire [63:0] R8972;
  wire [63:0] R8971;
  wire [63:0] R8970;
  wire [63:0] R8969;
  wire [63:0] R8968;
  wire [63:0] R8967;
  wire [63:0] R8966;
  wire [63:0] R8965;
  wire [63:0] R8964;
  wire [31:0] R8963;
  wire [63:0] R8962;
  wire [63:0] R8961;
  wire [63:0] R8960;
  wire [63:0] R8959;
  wire [63:0] R8958;
  wire [63:0] R8957;
  wire [31:0] R8956;
  wire [63:0] R8955;
  wire [63:0] R8954;
  wire [63:0] R8953;
  wire [63:0] R8952;
  wire [63:0] R8951;
  wire [63:0] R8950;
  wire [31:0] R8949;
  wire [63:0] R8948;
  wire [63:0] R8947;
  wire [63:0] R8946;
  wire [63:0] R8945;
  wire [63:0] R8944;
  wire [63:0] R8943;
  wire [31:0] R8942;
  wire [63:0] R8941;
  wire [63:0] R8940;
  wire [63:0] R8939;
  wire [63:0] R8938;
  wire [63:0] R8937;
  wire [63:0] R8936;
  wire [31:0] R8935;
  wire [63:0] R8934;
  wire [63:0] R8933;
  wire [63:0] R8932;
  wire [63:0] R8931;
  wire [63:0] R8930;
  wire [63:0] R8929;
  wire [31:0] R8928;
  wire [63:0] R8927;
  wire [63:0] R8926;
  wire [63:0] R8925;
  wire [63:0] R8924;
  wire [63:0] R8923;
  wire [63:0] R8922;
  wire [63:0] R8921;
  wire [63:0] R8920;
  wire [63:0] R8919;
  wire [63:0] R8918;
  wire [63:0] R8917;
  wire [63:0] R8916;
  wire [63:0] R8915;
  wire [63:0] R8914;
  wire [63:0] R8913;
  wire [63:0] R8912;
  wire [63:0] R8911;
  wire [63:0] R8910;
  wire [63:0] R8909;
  wire [63:0] R8908;
  wire [63:0] R8907;
  wire [31:0] R8906;
  wire [63:0] R8905;
  wire [63:0] R8904;
  wire [63:0] R8903;
  wire [63:0] R8902;
  wire [63:0] R8901;
  wire [63:0] R8900;
  wire [31:0] R8899;
  wire [63:0] R8898;
  wire [63:0] R8897;
  wire [63:0] R8896;
  wire [63:0] R8895;
  wire [63:0] R8894;
  wire [63:0] R8893;
  wire [31:0] R8892;
  wire [63:0] R8891;
  wire [63:0] R8890;
  wire [63:0] R8889;
  wire [63:0] R8888;
  wire [63:0] R8887;
  wire [63:0] R8886;
  wire [31:0] R8885;
  wire [63:0] R8884;
  wire [63:0] R8883;
  wire [63:0] R8882;
  wire [63:0] R8881;
  wire [63:0] R8880;
  wire [63:0] R8879;
  wire [31:0] R8878;
  wire [63:0] R8877;
  wire [63:0] R8876;
  wire [63:0] R8875;
  wire [63:0] R8874;
  wire [63:0] R8873;
  wire [63:0] R8872;
  wire [31:0] R8871;
  wire [63:0] R8870;
  wire [63:0] R8869;
  wire [63:0] R8868;
  wire [63:0] R8867;
  wire [63:0] R8866;
  wire [63:0] R8865;
  wire [31:0] R8864;
  wire [63:0] R8863;
  wire [63:0] R8862;
  wire [63:0] R8861;
  wire [63:0] R8860;
  wire [63:0] R8859;
  wire [63:0] R8858;
  wire [31:0] R8857;
  wire [63:0] R8856;
  wire [63:0] R8855;
  wire [63:0] R8854;
  wire [63:0] R8853;
  wire [63:0] R8852;
  wire [63:0] R8851;
  wire [31:0] R8850;
  wire [63:0] R8849;
  wire [63:0] R8848;
  wire [63:0] R8847;
  wire [63:0] R8846;
  wire [63:0] R8845;
  wire [63:0] R8844;
  wire [31:0] R8843;
  wire [31:0] R8842;
  wire [31:0] R8841;
  wire [63:0] R8840;
  wire [31:0] R8839;
  wire [31:0] R8838;
  wire [31:0] R8837;
  wire [63:0] R8836;
  wire [31:0] R8835;
  wire [31:0] R8834;
  wire [31:0] R8833;
  wire [63:0] R8832;
  wire [31:0] R8831;
  wire [31:0] R8830;
  wire [31:0] R8829;
  wire [63:0] R8828;
  wire [31:0] R8827;
  wire [31:0] R8826;
  wire [31:0] R8825;
  wire [63:0] R8824;
  wire [31:0] R8823;
  wire [31:0] R8822;
  wire [31:0] R8821;
  wire [63:0] R8820;
  wire [63:0] R8819;
  wire [63:0] R8818;
  wire [63:0] R8817;
  wire [63:0] R8816;
  wire [63:0] R8815;
  wire [63:0] R8814;
  wire [63:0] R8813;
  wire [63:0] R8812;
  wire [63:0] R8811;
  wire [63:0] R8810;
  wire [63:0] R8809;
  wire [63:0] R8808;
  wire [63:0] R8807;
  wire [63:0] R8806;
  wire [63:0] R8805;
  wire [63:0] R8804;
  wire [63:0] R8803;
  wire [63:0] R8802;
  wire [63:0] R8801;
  wire [63:0] R8800;
  wire [63:0] R8799;
  wire [63:0] R8798;
  wire [63:0] R8797;
  wire [63:0] R8796;
  wire [63:0] R8795;
  wire [63:0] R8794;
  wire [63:0] R8793;
  wire [63:0] R8792;
  wire [63:0] R8791;
  wire [63:0] R8790;
  wire [63:0] R8789;
  wire [63:0] R8788;
  wire [63:0] R8787;
  wire [63:0] R8786;
  wire [63:0] R8785;
  wire [63:0] R8784;
  wire [63:0] R8783;
  wire [63:0] R8782;
  wire [63:0] R8781;
  wire [63:0] R8780;
  wire [63:0] R8779;
  wire [63:0] R8778;
  wire [63:0] R8777;
  wire [63:0] R8776;
  wire [63:0] R8775;
  wire [63:0] R8774;
  wire [63:0] R8773;
  wire [63:0] R8772;
  wire [63:0] R8771;
  wire [63:0] R8770;
  wire [63:0] R8769;
  wire [31:0] R8768;
  wire [31:0] R8767;
  wire [31:0] R8766;
  wire [63:0] R8765;
  wire [31:0] R8764;
  wire [31:0] R8763;
  wire [31:0] R8762;
  wire [63:0] R8761;
  wire [31:0] R8760;
  wire [31:0] R8759;
  wire [31:0] R8758;
  wire [63:0] R8757;
  wire [31:0] R8756;
  wire [31:0] R8755;
  wire [31:0] R8754;
  wire [63:0] R8753;
  wire [31:0] R8752;
  wire [31:0] R8751;
  wire [31:0] R8750;
  wire [63:0] R8749;
  wire [31:0] R8748;
  wire [31:0] R8747;
  wire [31:0] R8746;
  wire [63:0] R8745;
  wire [31:0] R8744;
  wire [31:0] R8743;
  wire [31:0] R8742;
  wire [63:0] R8741;
  wire [31:0] R8740;
  wire [31:0] R8739;
  wire [31:0] R8738;
  wire [63:0] R8737;
  wire [31:0] R8736;
  wire [31:0] R8735;
  wire [31:0] R8734;
  wire [63:0] R8733;
  wire [63:0] R8732;
  wire [63:0] R8731;
  wire [63:0] R8730;
  wire [63:0] R8729;
  wire [63:0] R8728;
  wire [63:0] R8727;
  wire [63:0] R8726;
  wire [63:0] R8725;
  wire [63:0] R8724;
  wire [63:0] R8723;
  wire [63:0] R8722;
  wire [63:0] R8721;
  wire [63:0] R8720;
  wire [63:0] R8719;
  wire [63:0] R8718;
  wire [63:0] R8717;
  wire [63:0] R8716;
  wire [63:0] R8715;
  wire [63:0] R8714;
  wire [63:0] R8713;
  wire [63:0] R8712;
  wire [63:0] R8711;
  wire [63:0] R8710;
  wire [63:0] R8709;
  wire [63:0] R8708;
  wire [63:0] R8707;
  wire [63:0] R8706;
  wire [63:0] R8705;
  wire [63:0] R8704;
  wire [63:0] R8703;
  wire [63:0] R8702;
  wire [63:0] R8701;
  wire [63:0] R8700;
  wire [63:0] R8699;
  wire [63:0] R8698;
  wire [63:0] R8697;
  wire [63:0] R8696;
  wire [63:0] R8695;
  wire [63:0] R8694;
  wire [63:0] R8693;
  wire [63:0] R8692;
  wire [63:0] R8691;
  wire [63:0] R8690;
  wire [63:0] R8689;
  wire [63:0] R8688;
  wire [63:0] R8687;
  wire [63:0] R8686;
  wire [63:0] R8685;
  wire [63:0] R8684;
  wire [63:0] R8683;
  wire [63:0] R8682;
  wire [63:0] R8681;
  wire [63:0] R8680;
  wire [63:0] R8679;
  wire [63:0] R8678;
  wire [63:0] R8677;
  wire [63:0] R8676;
  wire [63:0] R8675;
  wire [63:0] R8674;
  wire [63:0] R8673;
  wire [63:0] R8672;
  wire [63:0] R8671;
  wire [63:0] R8670;
  wire [63:0] R8669;
  wire [63:0] R8668;
  wire [63:0] R8667;
  wire [63:0] R8666;
  wire [63:0] R8665;
  wire [63:0] R8664;
  wire [63:0] R8663;
  wire [63:0] R8662;
  wire [63:0] R8661;
  wire [63:0] R8660;
  wire [63:0] R8659;
  wire [63:0] R8658;
  wire [63:0] R8657;
  wire [63:0] R8656;
  wire [63:0] R8655;
  wire [63:0] R8654;
  wire [63:0] R8653;
  wire [63:0] R8652;
  wire [63:0] R8651;
  wire [63:0] R8650;
  wire [63:0] R8649;
  wire [63:0] R8648;
  wire [63:0] R8647;
  wire [63:0] R8646;
  wire [63:0] R8645;
  wire [63:0] R8644;
  wire [63:0] R8643;
  wire [63:0] R8642;
  wire [63:0] R8641;
  wire [63:0] R8640;
  wire [63:0] R8639;
  wire [63:0] R8638;
  wire [63:0] R8637;
  wire [63:0] R8636;
  wire [63:0] R8635;
  wire [63:0] R8634;
  wire [63:0] R8633;
  wire [63:0] R8632;
  wire [63:0] R8631;
  wire [63:0] R8630;
  wire [63:0] R8629;
  wire [63:0] R8628;
  wire [63:0] R8627;
  wire [63:0] R8626;
  wire [63:0] R8625;
  wire [63:0] R8624;
  wire [63:0] R8623;
  wire [63:0] R8622;
  wire [63:0] R8621;
  wire [63:0] R8620;
  wire [63:0] R8619;
  wire [63:0] R8618;
  wire [63:0] R8617;
  wire [63:0] R8616;
  wire [63:0] R8615;
  wire [63:0] R8614;
  wire [63:0] R8613;
  wire [63:0] R8612;
  wire [63:0] R8611;
  wire [63:0] R8610;
  wire [63:0] R8609;
  wire [63:0] R8608;
  wire [63:0] R8607;
  wire [63:0] R8606;
  wire [63:0] R8605;
  wire [63:0] R8604;
  wire [63:0] R8603;
  wire [63:0] R8602;
  wire [63:0] R8601;
  wire [63:0] R8600;
  wire [63:0] R8599;
  wire [63:0] R8598;
  wire [63:0] R8597;
  wire [63:0] R8596;
  wire [63:0] R8595;
  wire [63:0] R8594;
  wire [63:0] R8593;
  wire [63:0] R8592;
  wire [63:0] R8591;
  wire [63:0] R8590;
  wire [63:0] R8589;
  wire [63:0] R8588;
  wire [63:0] R8587;
  wire [63:0] R8586;
  wire [63:0] R8585;
  wire [63:0] R8584;
  wire [63:0] R8583;
  wire [63:0] R8582;
  wire [63:0] R8581;
  wire [63:0] R8580;
  wire [63:0] R8579;
  wire [63:0] R8578;
  wire [63:0] R8577;
  wire [63:0] R8576;
  wire [63:0] R8575;
  wire [63:0] R8574;
  wire [63:0] R8573;
  wire [63:0] R8572;
  wire [63:0] R8571;
  wire [63:0] R8570;
  wire [63:0] R8569;
  wire [63:0] R8568;
  wire [63:0] R8567;
  wire [63:0] R8566;
  wire [63:0] R8565;
  wire [63:0] R8564;
  wire [63:0] R8563;
  wire [63:0] R8562;
  wire [63:0] R8561;
  wire [63:0] R8560;
  wire [63:0] R8559;
  wire [63:0] R8558;
  wire [63:0] R8557;
  wire [63:0] R8556;
  wire [63:0] R8555;
  wire [63:0] R8554;
  wire [63:0] R8553;
  wire [63:0] R8552;
  wire [63:0] R8551;
  wire [63:0] R8550;
  wire [63:0] R8549;
  wire [63:0] R8548;
  wire [63:0] R8547;
  wire [63:0] R8546;
  wire [63:0] R8545;
  wire [63:0] R8544;
  wire [63:0] R8543;
  wire [63:0] R8542;
  wire [63:0] R8541;
  wire [63:0] R8540;
  wire [63:0] R8539;
  wire [63:0] R8538;
  wire [63:0] R8537;
  wire [63:0] R8536;
  wire [63:0] R8535;
  wire [63:0] R8534;
  wire [63:0] R8533;
  wire [63:0] R8532;
  wire [63:0] R8531;
  wire [63:0] R8530;
  wire [63:0] R8529;
  wire [63:0] R8528;
  wire [63:0] R8527;
  wire [63:0] R8526;
  wire [63:0] R8525;
  wire [63:0] R8524;
  wire [63:0] R8523;
  wire [63:0] R8522;
  wire [63:0] R8521;
  wire [63:0] R8520;
  wire [63:0] R8519;
  wire [63:0] R8518;
  wire [63:0] R8517;
  wire [63:0] R8516;
  wire [63:0] R8515;
  wire [63:0] R8514;
  wire [63:0] R8513;
  wire [63:0] R8512;
  wire [63:0] R8511;
  wire [63:0] R8510;
  wire [63:0] R8509;
  wire [63:0] R8508;
  wire [63:0] R8507;
  wire [63:0] R8506;
  wire [63:0] R8505;
  wire [63:0] R8504;
  wire [63:0] R8503;
  wire [63:0] R8502;
  wire [63:0] R8501;
  wire [63:0] R8500;
  wire [63:0] R8499;
  wire [63:0] R8498;
  wire [63:0] R8497;
  wire [63:0] R8496;
  wire [63:0] R8495;
  wire [63:0] R8494;
  wire [63:0] R8493;
  wire [63:0] R8492;
  wire [63:0] R8491;
  wire [63:0] R8490;
  wire [63:0] R8489;
  wire [63:0] R8488;
  wire [63:0] R8487;
  wire [63:0] R8486;
  wire [63:0] R8485;
  wire [63:0] R8484;
  wire [63:0] R8483;
  wire [63:0] R8482;
  wire [63:0] R8481;
  wire [63:0] R8480;
  wire [63:0] R8479;
  wire [63:0] R8478;
  wire [63:0] R8477;
  wire [63:0] R8476;
  wire [63:0] R8475;
  wire [63:0] R8474;
  wire [63:0] R8473;
  wire [63:0] R8472;
  wire [63:0] R8471;
  wire [63:0] R8470;
  wire [63:0] R8469;
  wire [63:0] R8468;
  wire [63:0] R8467;
  wire [63:0] R8466;
  wire [63:0] R8465;
  wire [63:0] R8464;
  wire [63:0] R8463;
  wire [63:0] R8462;
  wire [63:0] R8461;
  wire [63:0] R8460;
  wire [63:0] R8459;
  wire [63:0] R8458;
  wire [63:0] R8457;
  wire [63:0] R8456;
  wire [63:0] R8455;
  wire [63:0] R8454;
  wire [63:0] R8453;
  wire [63:0] R8452;
  wire [63:0] R8451;
  wire [63:0] R8450;
  wire [63:0] R8449;
  wire [63:0] R8448;
  wire [63:0] R8447;
  wire [63:0] R8446;
  wire [63:0] R8445;
  wire [63:0] R8444;
  wire [63:0] R8443;
  wire [63:0] R8442;
  wire [63:0] R8441;
  wire [63:0] R8440;
  wire [63:0] R8439;
  wire [0:0] R8438;
  wire [0:0] R8437;
  wire [0:0] R8436;
  wire [0:0] R8435;
  wire [0:0] R8434;
  wire [0:0] R8433;
  wire [0:0] R8432;
  wire [0:0] R8431;
  wire [0:0] R8430;
  wire [0:0] R8429;
  wire [0:0] R8428;
  wire [0:0] R8427;
  wire [0:0] R8426;
  wire [0:0] R8425;
  wire [0:0] R8424;
  wire [0:0] R8423;
  wire [0:0] R8422;
  wire [0:0] R8421;
  wire [0:0] R8420;
  wire [0:0] R8419;
  wire [0:0] R8418;
  wire [0:0] R8417;
  wire [0:0] R8416;
  wire [0:0] R8415;
  wire [0:0] R8414;
  wire [0:0] R8413;
  wire [0:0] R8412;
  wire [0:0] R8411;
  wire [0:0] R8410;
  wire [0:0] R8409;
  wire [0:0] R8408;
  wire [0:0] R8407;
  wire [0:0] R8406;
  wire [0:0] R8405;
  wire [0:0] R8404;
  wire [0:0] R8403;
  wire [0:0] R8402;
  wire [0:0] R8401;
  wire [0:0] R8400;
  wire [0:0] R8399;
  wire [0:0] R8398;
  wire [0:0] R8397;
  wire [0:0] R8396;
  wire [0:0] R8395;
  wire [0:0] R8394;
  wire [0:0] R8393;
  wire [0:0] R8392;
  wire [0:0] R8391;
  wire [0:0] R8390;
  wire [0:0] R8389;
  wire [0:0] R8388;
  wire [0:0] R8387;
  wire [0:0] R8386;
  wire [0:0] R8385;
  wire [0:0] R8384;
  wire [0:0] R8383;
  wire [0:0] R8382;
  wire [0:0] R8381;
  wire [0:0] R8380;
  wire [0:0] R8379;
  wire [0:0] R8378;
  wire [0:0] R8377;
  wire [0:0] R8376;
  wire [0:0] R8375;
  wire [0:0] R8374;
  wire [0:0] R8373;
  wire [63:0] R8372;
  wire [63:0] R8371;
  wire [63:0] R8370;
  wire [63:0] R8369;
  wire [63:0] R8368;
  wire [63:0] R8367;
  wire [63:0] R8366;
  wire [63:0] R8365;
  wire [63:0] R8364;
  wire [63:0] R8363;
  wire [63:0] R8362;
  wire [63:0] R8361;
  wire [63:0] R8360;
  wire [63:0] R8359;
  wire [63:0] R8358;
  wire [0:0] R8357;
  wire [0:0] R8356;
  wire [0:0] R8355;
  wire [0:0] R8354;
  wire [0:0] R8353;
  wire [0:0] R8352;
  wire [0:0] R8351;
  wire [0:0] R8350;
  wire [0:0] R8349;
  wire [0:0] R8348;
  wire [0:0] R8347;
  wire [0:0] R8346;
  wire [0:0] R8345;
  wire [0:0] R8344;
  wire [0:0] R8343;
  wire [0:0] R8342;
  wire [0:0] R8341;
  wire [0:0] R8340;
  wire [0:0] R8339;
  wire [0:0] R8338;
  wire [0:0] R8337;
  wire [0:0] R8336;
  wire [0:0] R8335;
  wire [0:0] R8334;
  wire [0:0] R8333;
  wire [0:0] R8332;
  wire [0:0] R8331;
  wire [0:0] R8330;
  wire [0:0] R8329;
  wire [0:0] R8328;
  wire [0:0] R8327;
  wire [0:0] R8326;
  wire [0:0] R8325;
  wire [0:0] R8324;
  wire [0:0] R8323;
  wire [0:0] R8322;
  wire [0:0] R8321;
  wire [0:0] R8320;
  wire [0:0] R8319;
  wire [0:0] R8318;
  wire [0:0] R8317;
  wire [0:0] R8316;
  wire [0:0] R8315;
  wire [0:0] R8314;
  wire [0:0] R8313;
  wire [0:0] R8312;
  wire [0:0] R8311;
  wire [0:0] R8310;
  wire [0:0] R8309;
  wire [0:0] R8308;
  wire [0:0] R8307;
  wire [0:0] R8306;
  wire [0:0] R8305;
  wire [0:0] R8304;
  wire [0:0] R8303;
  wire [0:0] R8302;
  wire [0:0] R8301;
  wire [0:0] R8300;
  wire [0:0] R8299;
  wire [0:0] R8298;
  wire [0:0] R8297;
  wire [0:0] R8296;
  wire [0:0] R8295;
  wire [0:0] R8294;
  wire [0:0] R8293;
  wire [0:0] R8292;
  wire [0:0] R8291;
  wire [0:0] R8290;
  wire [0:0] R8289;
  wire [0:0] R8288;
  wire [0:0] R8287;
  wire [0:0] R8286;
  wire [0:0] R8285;
  wire [0:0] R8284;
  wire [0:0] R8283;
  wire [0:0] R8282;
  wire [0:0] R8281;
  wire [0:0] R8280;
  wire [0:0] R8279;
  wire [0:0] R8278;
  wire [0:0] R8277;
  wire [0:0] R8276;
  wire [0:0] R8275;
  wire [0:0] R8274;
  wire [0:0] R8273;
  wire [0:0] R8272;
  wire [0:0] R8271;
  wire [0:0] R8270;
  wire [0:0] R8269;
  wire [0:0] R8268;
  wire [0:0] R8267;
  wire [0:0] R8266;
  wire [0:0] R8265;
  wire [0:0] R8264;
  wire [0:0] R8263;
  wire [0:0] R8262;
  wire [0:0] R8261;
  wire [0:0] R8260;
  wire [0:0] R8259;
  wire [63:0] R8258;
  wire [63:0] R8257;
  wire [63:0] R8256;
  wire [63:0] R8255;
  wire [63:0] R8254;
  wire [63:0] R8253;
  wire [63:0] R8252;
  wire [63:0] R8251;
  wire [63:0] R8250;
  wire [63:0] R8249;
  wire [63:0] R8248;
  wire [63:0] R8247;
  wire [63:0] R8246;
  wire [63:0] R8245;
  wire [63:0] R8244;
  wire [31:0] R8243;
  wire [31:0] R8242;
  wire [31:0] R8241;
  wire [31:0] R8240;
  wire [31:0] R8239;
  wire [63:0] R8238;
  wire [63:0] R8237;
  wire [63:0] R8236;
  wire [63:0] R8235;
  wire [63:0] R8234;
  wire [63:0] R8233;
  wire [63:0] R8232;
  wire [63:0] R8231;
  wire [63:0] R8230;
  wire [63:0] R8229;
  wire [63:0] R8228;
  wire [63:0] R8227;
  wire [63:0] R8226;
  wire [63:0] R8225;
  wire [63:0] R8224;
  wire [63:0] R8223;
  wire [63:0] R8222;
  wire [63:0] R8221;
  wire [63:0] R8220;
  wire [63:0] R8219;
  wire [63:0] R8218;
  wire [63:0] R8217;
  wire [63:0] R8216;
  wire [63:0] R8215;
  wire [63:0] R8214;
  wire [63:0] R8213;
  wire [63:0] R8212;
  wire [63:0] R8211;
  wire [63:0] R8210;
  wire [63:0] R8209;
  wire [63:0] R8208;
  wire [63:0] R8207;
  wire [63:0] R8206;
  wire [63:0] R8205;
  wire [63:0] R8204;
  wire [63:0] R8203;
  wire [63:0] R8202;
  wire [63:0] R8201;
  wire [63:0] R8200;
  wire [31:0] R8199;
  wire [31:0] R8198;
  wire [31:0] R8197;
  wire [31:0] R8196;
  wire [31:0] R8195;
  wire [31:0] R8194;
  wire [31:0] R8193;
  wire [31:0] R8192;
  wire [31:0] R8191;
  wire [31:0] R8190;
  wire [31:0] R8189;
  wire [31:0] R8188;
  wire [31:0] R8187;
  wire [31:0] R8186;
  wire [63:0] R8185;
  wire [31:0] R8184;
  wire [63:0] R8183;
  wire [63:0] R8182;
  wire [63:0] R8181;
  wire [63:0] R8180;
  wire [63:0] R8179;
  wire [63:0] R8178;
  wire [31:0] R8177;
  wire [63:0] R8176;
  wire [63:0] R8175;
  wire [63:0] R8174;
  wire [63:0] R8173;
  wire [63:0] R8172;
  wire [63:0] R8171;
  wire [63:0] R8170;
  wire [31:0] R8169;
  wire [31:0] R8168;
  wire [31:0] R8167;
  wire [63:0] R8166;
  wire [63:0] R8165;
  wire [63:0] R8164;
  wire [63:0] R8163;
  wire [63:0] R8162;
  wire [63:0] R8161;
  wire [63:0] R8160;
  wire [63:0] R8159;
  wire [63:0] R8158;
  wire [63:0] R8157;
  wire [63:0] R8156;
  wire [63:0] R8155;
  wire [63:0] R8154;
  wire [63:0] R8153;
  wire [63:0] R8152;
  wire [63:0] R8151;
  wire [63:0] R8150;
  wire [63:0] R8149;
  wire [63:0] R8148;
  wire [63:0] R8147;
  wire [63:0] R8146;
  wire [63:0] R8145;
  wire [63:0] R8144;
  wire [63:0] R8143;
  wire [0:0] R8142;
  wire [0:0] R8141;
  wire [0:0] R8140;
  wire [0:0] R8139;
  wire [0:0] R8138;
  wire [0:0] R8137;
  wire [0:0] R8136;
  wire [0:0] R8135;
  wire [0:0] R8134;
  wire [0:0] R8133;
  wire [0:0] R8132;
  wire [0:0] R8131;
  wire [0:0] R8130;
  wire [0:0] R8129;
  wire [0:0] R8128;
  wire [0:0] R8127;
  wire [0:0] R8126;
  wire [0:0] R8125;
  wire [0:0] R8124;
  wire [0:0] R8123;
  wire [0:0] R8122;
  wire [0:0] R8121;
  wire [0:0] R8120;
  wire [0:0] R8119;
  wire [0:0] R8118;
  wire [63:0] R8117;
  wire [31:0] R8116;
  wire [31:0] R8115;
  wire [31:0] R8114;
  wire [31:0] R8113;
  wire [31:0] R8112;
  wire [31:0] R8111;
  wire [31:0] R8110;
  wire [31:0] R8109;
  wire [31:0] R8108;
  wire [31:0] R8107;
  wire [31:0] R8106;
  wire [31:0] R8105;
  wire [31:0] R8104;
  wire [31:0] R8103;
  wire [31:0] R8102;
  wire [31:0] R8101;
  wire [31:0] R8100;
  wire [31:0] R8099;
  wire [31:0] R8098;
  wire [63:0] R8097;
  wire [63:0] R8096;
  wire [63:0] R8095;
  wire [31:0] R8094;
  wire [31:0] R8093;
  wire [31:0] R8092;
  wire [31:0] R8091;
  wire [31:0] R8090;
  wire [31:0] R8089;
  wire [31:0] R8088;
  wire [31:0] R8087;
  wire [31:0] R8086;
  wire [31:0] R8085;
  wire [31:0] R8084;
  wire [31:0] R8083;
  wire [31:0] R8082;
  wire [31:0] R8081;
  wire [31:0] R8080;
  wire [31:0] R8079;
  wire [31:0] R8078;
  wire [31:0] R8077;
  wire [31:0] R8076;
  wire [31:0] R8075;
  wire [31:0] R8074;
  wire [31:0] R8073;
  wire [31:0] R8072;
  wire [31:0] R8071;
  wire [31:0] R8070;
  wire [31:0] R8069;
  wire [63:0] R8068;
  wire [31:0] R8067;
  wire [31:0] R8066;
  wire [63:0] R8065;
  wire [31:0] R8064;
  wire [63:0] R8063;
  wire [63:0] R8062;
  wire [63:0] R8061;
  wire [63:0] R8060;
  wire [63:0] R8059;
  wire [63:0] R8058;
  wire [31:0] R8057;
  wire [63:0] R8056;
  wire [63:0] R8055;
  wire [63:0] R8054;
  wire [63:0] R8053;
  wire [63:0] R8052;
  wire [63:0] R8051;
  wire [63:0] R8050;
  wire [31:0] R8049;
  wire [31:0] R8048;
  wire [31:0] R8047;
  wire [63:0] R8046;
  wire [63:0] R8045;
  wire [63:0] R8044;
  wire [63:0] R8043;
  wire [63:0] R8042;
  wire [63:0] R8041;
  wire [63:0] R8040;
  wire [63:0] R8039;
  wire [63:0] R8038;
  wire [63:0] R8037;
  wire [63:0] R8036;
  wire [63:0] R8035;
  wire [63:0] R8034;
  wire [63:0] R8033;
  wire [63:0] R8032;
  wire [63:0] R8031;
  wire [63:0] R8030;
  wire [63:0] R8029;
  wire [63:0] R8028;
  wire [63:0] R8027;
  wire [63:0] R8026;
  wire [63:0] R8025;
  wire [63:0] R8024;
  wire [63:0] R8023;
  wire [0:0] R8022;
  wire [0:0] R8021;
  wire [0:0] R8020;
  wire [0:0] R8019;
  wire [0:0] R8018;
  wire [0:0] R8017;
  wire [0:0] R8016;
  wire [0:0] R8015;
  wire [0:0] R8014;
  wire [0:0] R8013;
  wire [0:0] R8012;
  wire [0:0] R8011;
  wire [0:0] R8010;
  wire [0:0] R8009;
  wire [0:0] R8008;
  wire [0:0] R8007;
  wire [0:0] R8006;
  wire [0:0] R8005;
  wire [0:0] R8004;
  wire [0:0] R8003;
  wire [0:0] R8002;
  wire [0:0] R8001;
  wire [0:0] R8000;
  wire [0:0] R7999;
  wire [0:0] R7998;
  wire [0:0] R7997;
  wire [0:0] R7996;
  wire [0:0] R7995;
  wire [0:0] R7994;
  wire [0:0] R7993;
  wire [0:0] R7992;
  wire [0:0] R7991;
  wire [0:0] R7990;
  wire [0:0] R7989;
  wire [0:0] R7988;
  wire [0:0] R7987;
  wire [0:0] R7986;
  wire [0:0] R7985;
  wire [0:0] R7984;
  wire [63:0] R7983;
  wire [31:0] R7982;
  wire [31:0] R7981;
  wire [31:0] R7980;
  wire [31:0] R7979;
  wire [31:0] R7978;
  wire [31:0] R7977;
  wire [31:0] R7976;
  wire [31:0] R7975;
  wire [31:0] R7974;
  wire [31:0] R7973;
  wire [31:0] R7972;
  wire [31:0] R7971;
  wire [31:0] R7970;
  wire [31:0] R7969;
  wire [31:0] R7968;
  wire [31:0] R7967;
  wire [31:0] R7966;
  wire [31:0] R7965;
  wire [31:0] R7964;
  wire [31:0] R7963;
  wire [31:0] R7962;
  wire [31:0] R7961;
  wire [31:0] R7960;
  wire [31:0] R7959;
  wire [31:0] R7958;
  wire [31:0] R7957;
  wire [31:0] R7956;
  wire [31:0] R7955;
  wire [31:0] R7954;
  wire [31:0] R7953;
  wire [31:0] R7952;
  wire [31:0] R7951;
  wire [31:0] R7950;
  wire [63:0] R7949;
  wire [63:0] R7948;
  wire [63:0] R7947;
  wire [31:0] R7946;
  wire [31:0] R7945;
  wire [31:0] R7944;
  wire [31:0] R7943;
  wire [31:0] R7942;
  wire [31:0] R7941;
  wire [31:0] R7940;
  wire [31:0] R7939;
  wire [31:0] R7938;
  wire [31:0] R7937;
  wire [31:0] R7936;
  wire [31:0] R7935;
  wire [31:0] R7934;
  wire [31:0] R7933;
  wire [31:0] R7932;
  wire [31:0] R7931;
  wire [31:0] R7930;
  wire [31:0] R7929;
  wire [31:0] R7928;
  wire [31:0] R7927;
  wire [31:0] R7926;
  wire [31:0] R7925;
  wire [31:0] R7924;
  wire [31:0] R7923;
  wire [31:0] R7922;
  wire [31:0] R7921;
  wire [31:0] R7920;
  wire [31:0] R7919;
  wire [31:0] R7918;
  wire [31:0] R7917;
  wire [31:0] R7916;
  wire [31:0] R7915;
  wire [31:0] R7914;
  wire [31:0] R7913;
  wire [31:0] R7912;
  wire [31:0] R7911;
  wire [31:0] R7910;
  wire [31:0] R7909;
  wire [31:0] R7908;
  wire [31:0] R7907;
  wire [63:0] R7906;
  wire [31:0] R7905;
  wire [31:0] R7904;
  wire [63:0] R7903;
  wire [31:0] R7902;
  wire [63:0] R7901;
  wire [63:0] R7900;
  wire [63:0] R7899;
  wire [63:0] R7898;
  wire [63:0] R7897;
  wire [63:0] R7896;
  wire [31:0] R7895;
  wire [63:0] R7894;
  wire [63:0] R7893;
  wire [63:0] R7892;
  wire [63:0] R7891;
  wire [63:0] R7890;
  wire [63:0] R7889;
  wire [63:0] R7888;
  wire [31:0] R7887;
  wire [31:0] R7886;
  wire [31:0] R7885;
  wire [63:0] R7884;
  wire [63:0] R7883;
  wire [63:0] R7882;
  wire [63:0] R7881;
  wire [63:0] R7880;
  wire [63:0] R7879;
  wire [63:0] R7878;
  wire [63:0] R7877;
  wire [63:0] R7876;
  wire [63:0] R7875;
  wire [63:0] R7874;
  wire [63:0] R7873;
  wire [63:0] R7872;
  wire [63:0] R7871;
  wire [63:0] R7870;
  wire [63:0] R7869;
  wire [63:0] R7868;
  wire [63:0] R7867;
  wire [63:0] R7866;
  wire [63:0] R7865;
  wire [63:0] R7864;
  wire [63:0] R7863;
  wire [63:0] R7862;
  wire [63:0] R7861;
  wire [0:0] R7860;
  wire [0:0] R7859;
  wire [0:0] R7858;
  wire [0:0] R7857;
  wire [0:0] R7856;
  wire [0:0] R7855;
  wire [0:0] R7854;
  wire [0:0] R7853;
  wire [0:0] R7852;
  wire [0:0] R7851;
  wire [0:0] R7850;
  wire [0:0] R7849;
  wire [0:0] R7848;
  wire [0:0] R7847;
  wire [0:0] R7846;
  wire [0:0] R7845;
  wire [0:0] R7844;
  wire [0:0] R7843;
  wire [0:0] R7842;
  wire [0:0] R7841;
  wire [0:0] R7840;
  wire [0:0] R7839;
  wire [0:0] R7838;
  wire [0:0] R7837;
  wire [0:0] R7836;
  wire [0:0] R7835;
  wire [0:0] R7834;
  wire [0:0] R7833;
  wire [0:0] R7832;
  wire [0:0] R7831;
  wire [0:0] R7830;
  wire [0:0] R7829;
  wire [0:0] R7828;
  wire [0:0] R7827;
  wire [0:0] R7826;
  wire [0:0] R7825;
  wire [0:0] R7824;
  wire [0:0] R7823;
  wire [0:0] R7822;
  wire [0:0] R7821;
  wire [0:0] R7820;
  wire [0:0] R7819;
  wire [0:0] R7818;
  wire [0:0] R7817;
  wire [0:0] R7816;
  wire [0:0] R7815;
  wire [0:0] R7814;
  wire [0:0] R7813;
  wire [0:0] R7812;
  wire [0:0] R7811;
  wire [0:0] R7810;
  wire [0:0] R7809;
  wire [0:0] R7808;
  wire [63:0] R7807;
  wire [31:0] R7806;
  wire [31:0] R7805;
  wire [31:0] R7804;
  wire [31:0] R7803;
  wire [31:0] R7802;
  wire [31:0] R7801;
  wire [31:0] R7800;
  wire [31:0] R7799;
  wire [31:0] R7798;
  wire [31:0] R7797;
  wire [31:0] R7796;
  wire [31:0] R7795;
  wire [31:0] R7794;
  wire [31:0] R7793;
  wire [31:0] R7792;
  wire [31:0] R7791;
  wire [31:0] R7790;
  wire [31:0] R7789;
  wire [31:0] R7788;
  wire [31:0] R7787;
  wire [31:0] R7786;
  wire [31:0] R7785;
  wire [31:0] R7784;
  wire [31:0] R7783;
  wire [31:0] R7782;
  wire [31:0] R7781;
  wire [31:0] R7780;
  wire [31:0] R7779;
  wire [31:0] R7778;
  wire [31:0] R7777;
  wire [31:0] R7776;
  wire [31:0] R7775;
  wire [31:0] R7774;
  wire [31:0] R7773;
  wire [31:0] R7772;
  wire [31:0] R7771;
  wire [31:0] R7770;
  wire [31:0] R7769;
  wire [31:0] R7768;
  wire [31:0] R7767;
  wire [31:0] R7766;
  wire [31:0] R7765;
  wire [31:0] R7764;
  wire [31:0] R7763;
  wire [31:0] R7762;
  wire [31:0] R7761;
  wire [31:0] R7760;
  wire [63:0] R7759;
  wire [63:0] R7758;
  wire [63:0] R7757;
  wire [31:0] R7756;
  wire [31:0] R7755;
  wire [31:0] R7754;
  wire [31:0] R7753;
  wire [31:0] R7752;
  wire [31:0] R7751;
  wire [31:0] R7750;
  wire [31:0] R7749;
  wire [31:0] R7748;
  wire [31:0] R7747;
  wire [31:0] R7746;
  wire [31:0] R7745;
  wire [31:0] R7744;
  wire [31:0] R7743;
  wire [31:0] R7742;
  wire [31:0] R7741;
  wire [31:0] R7740;
  wire [31:0] R7739;
  wire [31:0] R7738;
  wire [31:0] R7737;
  wire [31:0] R7736;
  wire [31:0] R7735;
  wire [31:0] R7734;
  wire [31:0] R7733;
  wire [31:0] R7732;
  wire [31:0] R7731;
  wire [31:0] R7730;
  wire [31:0] R7729;
  wire [31:0] R7728;
  wire [31:0] R7727;
  wire [31:0] R7726;
  wire [31:0] R7725;
  wire [31:0] R7724;
  wire [31:0] R7723;
  wire [31:0] R7722;
  wire [31:0] R7721;
  wire [31:0] R7720;
  wire [31:0] R7719;
  wire [31:0] R7718;
  wire [31:0] R7717;
  wire [31:0] R7716;
  wire [31:0] R7715;
  wire [31:0] R7714;
  wire [31:0] R7713;
  wire [31:0] R7712;
  wire [31:0] R7711;
  wire [31:0] R7710;
  wire [31:0] R7709;
  wire [31:0] R7708;
  wire [31:0] R7707;
  wire [31:0] R7706;
  wire [31:0] R7705;
  wire [31:0] R7704;
  wire [31:0] R7703;
  wire [63:0] R7702;
  wire [31:0] R7701;
  wire [31:0] R7700;
  wire [63:0] R7699;
  wire [31:0] R7698;
  wire [63:0] R7697;
  wire [63:0] R7696;
  wire [63:0] R7695;
  wire [63:0] R7694;
  wire [63:0] R7693;
  wire [63:0] R7692;
  wire [31:0] R7691;
  wire [63:0] R7690;
  wire [63:0] R7689;
  wire [63:0] R7688;
  wire [63:0] R7687;
  wire [63:0] R7686;
  wire [63:0] R7685;
  wire [63:0] R7684;
  wire [31:0] R7683;
  wire [31:0] R7682;
  wire [31:0] R7681;
  wire [63:0] R7680;
  wire [63:0] R7679;
  wire [63:0] R7678;
  wire [63:0] R7677;
  wire [63:0] R7676;
  wire [63:0] R7675;
  wire [63:0] R7674;
  wire [63:0] R7673;
  wire [63:0] R7672;
  wire [63:0] R7671;
  wire [63:0] R7670;
  wire [63:0] R7669;
  wire [63:0] R7668;
  wire [63:0] R7667;
  wire [63:0] R7666;
  wire [63:0] R7665;
  wire [63:0] R7664;
  wire [63:0] R7663;
  wire [63:0] R7662;
  wire [63:0] R7661;
  wire [63:0] R7660;
  wire [63:0] R7659;
  wire [63:0] R7658;
  wire [63:0] R7657;
  wire [0:0] R7656;
  wire [0:0] R7655;
  wire [0:0] R7654;
  wire [0:0] R7653;
  wire [0:0] R7652;
  wire [0:0] R7651;
  wire [0:0] R7650;
  wire [0:0] R7649;
  wire [0:0] R7648;
  wire [0:0] R7647;
  wire [0:0] R7646;
  wire [0:0] R7645;
  wire [0:0] R7644;
  wire [0:0] R7643;
  wire [0:0] R7642;
  wire [0:0] R7641;
  wire [0:0] R7640;
  wire [0:0] R7639;
  wire [0:0] R7638;
  wire [0:0] R7637;
  wire [0:0] R7636;
  wire [0:0] R7635;
  wire [0:0] R7634;
  wire [0:0] R7633;
  wire [0:0] R7632;
  wire [0:0] R7631;
  wire [0:0] R7630;
  wire [0:0] R7629;
  wire [0:0] R7628;
  wire [0:0] R7627;
  wire [0:0] R7626;
  wire [0:0] R7625;
  wire [0:0] R7624;
  wire [0:0] R7623;
  wire [0:0] R7622;
  wire [0:0] R7621;
  wire [0:0] R7620;
  wire [0:0] R7619;
  wire [0:0] R7618;
  wire [0:0] R7617;
  wire [0:0] R7616;
  wire [0:0] R7615;
  wire [0:0] R7614;
  wire [0:0] R7613;
  wire [0:0] R7612;
  wire [0:0] R7611;
  wire [0:0] R7610;
  wire [0:0] R7609;
  wire [0:0] R7608;
  wire [0:0] R7607;
  wire [0:0] R7606;
  wire [0:0] R7605;
  wire [0:0] R7604;
  wire [0:0] R7603;
  wire [0:0] R7602;
  wire [0:0] R7601;
  wire [0:0] R7600;
  wire [0:0] R7599;
  wire [0:0] R7598;
  wire [0:0] R7597;
  wire [0:0] R7596;
  wire [0:0] R7595;
  wire [0:0] R7594;
  wire [0:0] R7593;
  wire [0:0] R7592;
  wire [0:0] R7591;
  wire [0:0] R7590;
  wire [63:0] R7589;
  wire [31:0] R7588;
  wire [31:0] R7587;
  wire [31:0] R7586;
  wire [31:0] R7585;
  wire [31:0] R7584;
  wire [31:0] R7583;
  wire [31:0] R7582;
  wire [31:0] R7581;
  wire [31:0] R7580;
  wire [31:0] R7579;
  wire [31:0] R7578;
  wire [31:0] R7577;
  wire [31:0] R7576;
  wire [31:0] R7575;
  wire [31:0] R7574;
  wire [31:0] R7573;
  wire [31:0] R7572;
  wire [31:0] R7571;
  wire [31:0] R7570;
  wire [31:0] R7569;
  wire [31:0] R7568;
  wire [31:0] R7567;
  wire [31:0] R7566;
  wire [31:0] R7565;
  wire [31:0] R7564;
  wire [31:0] R7563;
  wire [31:0] R7562;
  wire [31:0] R7561;
  wire [31:0] R7560;
  wire [31:0] R7559;
  wire [31:0] R7558;
  wire [31:0] R7557;
  wire [31:0] R7556;
  wire [31:0] R7555;
  wire [31:0] R7554;
  wire [31:0] R7553;
  wire [31:0] R7552;
  wire [31:0] R7551;
  wire [31:0] R7550;
  wire [31:0] R7549;
  wire [31:0] R7548;
  wire [31:0] R7547;
  wire [31:0] R7546;
  wire [31:0] R7545;
  wire [31:0] R7544;
  wire [31:0] R7543;
  wire [31:0] R7542;
  wire [31:0] R7541;
  wire [31:0] R7540;
  wire [31:0] R7539;
  wire [31:0] R7538;
  wire [31:0] R7537;
  wire [31:0] R7536;
  wire [31:0] R7535;
  wire [31:0] R7534;
  wire [31:0] R7533;
  wire [31:0] R7532;
  wire [31:0] R7531;
  wire [31:0] R7530;
  wire [31:0] R7529;
  wire [31:0] R7528;
  wire [63:0] R7527;
  wire [63:0] R7526;
  wire [63:0] R7525;
  wire [31:0] R7524;
  wire [31:0] R7523;
  wire [31:0] R7522;
  wire [31:0] R7521;
  wire [31:0] R7520;
  wire [31:0] R7519;
  wire [31:0] R7518;
  wire [31:0] R7517;
  wire [31:0] R7516;
  wire [31:0] R7515;
  wire [31:0] R7514;
  wire [31:0] R7513;
  wire [31:0] R7512;
  wire [31:0] R7511;
  wire [31:0] R7510;
  wire [31:0] R7509;
  wire [31:0] R7508;
  wire [31:0] R7507;
  wire [31:0] R7506;
  wire [31:0] R7505;
  wire [31:0] R7504;
  wire [31:0] R7503;
  wire [31:0] R7502;
  wire [31:0] R7501;
  wire [31:0] R7500;
  wire [31:0] R7499;
  wire [31:0] R7498;
  wire [31:0] R7497;
  wire [31:0] R7496;
  wire [31:0] R7495;
  wire [31:0] R7494;
  wire [31:0] R7493;
  wire [31:0] R7492;
  wire [31:0] R7491;
  wire [31:0] R7490;
  wire [31:0] R7489;
  wire [31:0] R7488;
  wire [31:0] R7487;
  wire [31:0] R7486;
  wire [31:0] R7485;
  wire [31:0] R7484;
  wire [31:0] R7483;
  wire [31:0] R7482;
  wire [31:0] R7481;
  wire [31:0] R7480;
  wire [31:0] R7479;
  wire [31:0] R7478;
  wire [31:0] R7477;
  wire [31:0] R7476;
  wire [31:0] R7475;
  wire [31:0] R7474;
  wire [31:0] R7473;
  wire [31:0] R7472;
  wire [31:0] R7471;
  wire [31:0] R7470;
  wire [31:0] R7469;
  wire [31:0] R7468;
  wire [31:0] R7467;
  wire [31:0] R7466;
  wire [31:0] R7465;
  wire [31:0] R7464;
  wire [31:0] R7463;
  wire [31:0] R7462;
  wire [31:0] R7461;
  wire [31:0] R7460;
  wire [31:0] R7459;
  wire [31:0] R7458;
  wire [31:0] R7457;
  wire [63:0] R7456;
  wire [31:0] R7455;
  wire [31:0] R7454;
  wire [63:0] R7453;
  wire [31:0] R7452;
  wire [63:0] R7451;
  wire [63:0] R7450;
  wire [63:0] R7449;
  wire [63:0] R7448;
  wire [63:0] R7447;
  wire [63:0] R7446;
  wire [31:0] R7445;
  wire [63:0] R7444;
  wire [63:0] R7443;
  wire [63:0] R7442;
  wire [63:0] R7441;
  wire [63:0] R7440;
  wire [63:0] R7439;
  wire [63:0] R7438;
  wire [31:0] R7437;
  wire [31:0] R7436;
  wire [31:0] R7435;
  wire [63:0] R7434;
  wire [63:0] R7433;
  wire [63:0] R7432;
  wire [63:0] R7431;
  wire [63:0] R7430;
  wire [63:0] R7429;
  wire [63:0] R7428;
  wire [63:0] R7427;
  wire [63:0] R7426;
  wire [63:0] R7425;
  wire [63:0] R7424;
  wire [63:0] R7423;
  wire [63:0] R7422;
  wire [63:0] R7421;
  wire [63:0] R7420;
  wire [63:0] R7419;
  wire [63:0] R7418;
  wire [63:0] R7417;
  wire [63:0] R7416;
  wire [63:0] R7415;
  wire [63:0] R7414;
  wire [63:0] R7413;
  wire [63:0] R7412;
  wire [63:0] R7411;
  wire [0:0] R7410;
  wire [0:0] R7409;
  wire [0:0] R7408;
  wire [0:0] R7407;
  wire [0:0] R7406;
  wire [0:0] R7405;
  wire [0:0] R7404;
  wire [0:0] R7403;
  wire [0:0] R7402;
  wire [0:0] R7401;
  wire [0:0] R7400;
  wire [0:0] R7399;
  wire [0:0] R7398;
  wire [0:0] R7397;
  wire [0:0] R7396;
  wire [0:0] R7395;
  wire [0:0] R7394;
  wire [0:0] R7393;
  wire [0:0] R7392;
  wire [0:0] R7391;
  wire [0:0] R7390;
  wire [0:0] R7389;
  wire [0:0] R7388;
  wire [0:0] R7387;
  wire [0:0] R7386;
  wire [0:0] R7385;
  wire [0:0] R7384;
  wire [0:0] R7383;
  wire [0:0] R7382;
  wire [0:0] R7381;
  wire [0:0] R7380;
  wire [0:0] R7379;
  wire [0:0] R7378;
  wire [0:0] R7377;
  wire [0:0] R7376;
  wire [0:0] R7375;
  wire [0:0] R7374;
  wire [0:0] R7373;
  wire [0:0] R7372;
  wire [0:0] R7371;
  wire [0:0] R7370;
  wire [0:0] R7369;
  wire [0:0] R7368;
  wire [0:0] R7367;
  wire [0:0] R7366;
  wire [0:0] R7365;
  wire [0:0] R7364;
  wire [0:0] R7363;
  wire [0:0] R7362;
  wire [0:0] R7361;
  wire [0:0] R7360;
  wire [0:0] R7359;
  wire [0:0] R7358;
  wire [0:0] R7357;
  wire [0:0] R7356;
  wire [0:0] R7355;
  wire [0:0] R7354;
  wire [0:0] R7353;
  wire [0:0] R7352;
  wire [0:0] R7351;
  wire [0:0] R7350;
  wire [0:0] R7349;
  wire [0:0] R7348;
  wire [0:0] R7347;
  wire [0:0] R7346;
  wire [0:0] R7345;
  wire [0:0] R7344;
  wire [0:0] R7343;
  wire [0:0] R7342;
  wire [0:0] R7341;
  wire [0:0] R7340;
  wire [0:0] R7339;
  wire [0:0] R7338;
  wire [0:0] R7337;
  wire [0:0] R7336;
  wire [0:0] R7335;
  wire [0:0] R7334;
  wire [0:0] R7333;
  wire [0:0] R7332;
  wire [0:0] R7331;
  wire [0:0] R7330;
  wire [63:0] R7329;
  wire [31:0] R7328;
  wire [31:0] R7327;
  wire [31:0] R7326;
  wire [31:0] R7325;
  wire [31:0] R7324;
  wire [31:0] R7323;
  wire [31:0] R7322;
  wire [31:0] R7321;
  wire [31:0] R7320;
  wire [31:0] R7319;
  wire [31:0] R7318;
  wire [31:0] R7317;
  wire [31:0] R7316;
  wire [31:0] R7315;
  wire [31:0] R7314;
  wire [31:0] R7313;
  wire [31:0] R7312;
  wire [31:0] R7311;
  wire [31:0] R7310;
  wire [31:0] R7309;
  wire [31:0] R7308;
  wire [31:0] R7307;
  wire [31:0] R7306;
  wire [31:0] R7305;
  wire [31:0] R7304;
  wire [31:0] R7303;
  wire [31:0] R7302;
  wire [31:0] R7301;
  wire [31:0] R7300;
  wire [31:0] R7299;
  wire [31:0] R7298;
  wire [31:0] R7297;
  wire [31:0] R7296;
  wire [31:0] R7295;
  wire [31:0] R7294;
  wire [31:0] R7293;
  wire [31:0] R7292;
  wire [31:0] R7291;
  wire [31:0] R7290;
  wire [31:0] R7289;
  wire [31:0] R7288;
  wire [31:0] R7287;
  wire [31:0] R7286;
  wire [31:0] R7285;
  wire [31:0] R7284;
  wire [31:0] R7283;
  wire [31:0] R7282;
  wire [31:0] R7281;
  wire [31:0] R7280;
  wire [31:0] R7279;
  wire [31:0] R7278;
  wire [31:0] R7277;
  wire [31:0] R7276;
  wire [31:0] R7275;
  wire [31:0] R7274;
  wire [31:0] R7273;
  wire [31:0] R7272;
  wire [31:0] R7271;
  wire [31:0] R7270;
  wire [31:0] R7269;
  wire [31:0] R7268;
  wire [31:0] R7267;
  wire [31:0] R7266;
  wire [31:0] R7265;
  wire [31:0] R7264;
  wire [31:0] R7263;
  wire [31:0] R7262;
  wire [31:0] R7261;
  wire [31:0] R7260;
  wire [31:0] R7259;
  wire [31:0] R7258;
  wire [31:0] R7257;
  wire [31:0] R7256;
  wire [31:0] R7255;
  wire [31:0] R7254;
  wire [63:0] R7253;
  wire [63:0] R7252;
  wire [63:0] R7251;
  wire [31:0] R7250;
  wire [31:0] R7249;
  wire [31:0] R7248;
  wire [31:0] R7247;
  wire [31:0] R7246;
  wire [31:0] R7245;
  wire [31:0] R7244;
  wire [31:0] R7243;
  wire [31:0] R7242;
  wire [31:0] R7241;
  wire [31:0] R7240;
  wire [31:0] R7239;
  wire [31:0] R7238;
  wire [31:0] R7237;
  wire [31:0] R7236;
  wire [31:0] R7235;
  wire [31:0] R7234;
  wire [31:0] R7233;
  wire [31:0] R7232;
  wire [31:0] R7231;
  wire [31:0] R7230;
  wire [31:0] R7229;
  wire [31:0] R7228;
  wire [31:0] R7227;
  wire [31:0] R7226;
  wire [31:0] R7225;
  wire [31:0] R7224;
  wire [31:0] R7223;
  wire [31:0] R7222;
  wire [31:0] R7221;
  wire [31:0] R7220;
  wire [31:0] R7219;
  wire [31:0] R7218;
  wire [31:0] R7217;
  wire [31:0] R7216;
  wire [31:0] R7215;
  wire [31:0] R7214;
  wire [31:0] R7213;
  wire [31:0] R7212;
  wire [31:0] R7211;
  wire [31:0] R7210;
  wire [31:0] R7209;
  wire [31:0] R7208;
  wire [31:0] R7207;
  wire [31:0] R7206;
  wire [31:0] R7205;
  wire [31:0] R7204;
  wire [31:0] R7203;
  wire [31:0] R7202;
  wire [31:0] R7201;
  wire [31:0] R7200;
  wire [31:0] R7199;
  wire [31:0] R7198;
  wire [31:0] R7197;
  wire [31:0] R7196;
  wire [31:0] R7195;
  wire [31:0] R7194;
  wire [31:0] R7193;
  wire [31:0] R7192;
  wire [31:0] R7191;
  wire [31:0] R7190;
  wire [31:0] R7189;
  wire [31:0] R7188;
  wire [31:0] R7187;
  wire [31:0] R7186;
  wire [31:0] R7185;
  wire [31:0] R7184;
  wire [31:0] R7183;
  wire [31:0] R7182;
  wire [31:0] R7181;
  wire [31:0] R7180;
  wire [31:0] R7179;
  wire [31:0] R7178;
  wire [31:0] R7177;
  wire [31:0] R7176;
  wire [31:0] R7175;
  wire [31:0] R7174;
  wire [31:0] R7173;
  wire [31:0] R7172;
  wire [31:0] R7171;
  wire [31:0] R7170;
  wire [31:0] R7169;
  wire [63:0] R7168;
  wire [31:0] R7167;
  wire [31:0] R7166;
  wire [63:0] R7165;
  wire [31:0] R7164;
  wire [63:0] R7163;
  wire [63:0] R7162;
  wire [63:0] R7161;
  wire [63:0] R7160;
  wire [63:0] R7159;
  wire [63:0] R7158;
  wire [31:0] R7157;
  wire [63:0] R7156;
  wire [63:0] R7155;
  wire [63:0] R7154;
  wire [63:0] R7153;
  wire [63:0] R7152;
  wire [63:0] R7151;
  wire [63:0] R7150;
  wire [31:0] R7149;
  wire [31:0] R7148;
  wire [31:0] R7147;
  wire [63:0] R7146;
  wire [63:0] R7145;
  wire [63:0] R7144;
  wire [63:0] R7143;
  wire [63:0] R7142;
  wire [63:0] R7141;
  wire [63:0] R7140;
  wire [63:0] R7139;
  wire [63:0] R7138;
  wire [63:0] R7137;
  wire [63:0] R7136;
  wire [63:0] R7135;
  wire [63:0] R7134;
  wire [63:0] R7133;
  wire [63:0] R7132;
  wire [63:0] R7131;
  wire [63:0] R7130;
  wire [63:0] R7129;
  wire [63:0] R7128;
  wire [63:0] R7127;
  wire [63:0] R7126;
  wire [63:0] R7125;
  wire [63:0] R7124;
  wire [63:0] R7123;
  wire [0:0] R7122;
  wire [0:0] R7121;
  wire [0:0] R7120;
  wire [0:0] R7119;
  wire [0:0] R7118;
  wire [0:0] R7117;
  wire [0:0] R7116;
  wire [0:0] R7115;
  wire [0:0] R7114;
  wire [0:0] R7113;
  wire [0:0] R7112;
  wire [0:0] R7111;
  wire [0:0] R7110;
  wire [0:0] R7109;
  wire [0:0] R7108;
  wire [0:0] R7107;
  wire [0:0] R7106;
  wire [0:0] R7105;
  wire [0:0] R7104;
  wire [0:0] R7103;
  wire [0:0] R7102;
  wire [0:0] R7101;
  wire [0:0] R7100;
  wire [0:0] R7099;
  wire [0:0] R7098;
  wire [0:0] R7097;
  wire [0:0] R7096;
  wire [0:0] R7095;
  wire [0:0] R7094;
  wire [0:0] R7093;
  wire [0:0] R7092;
  wire [0:0] R7091;
  wire [0:0] R7090;
  wire [0:0] R7089;
  wire [0:0] R7088;
  wire [0:0] R7087;
  wire [0:0] R7086;
  wire [0:0] R7085;
  wire [0:0] R7084;
  wire [0:0] R7083;
  wire [0:0] R7082;
  wire [0:0] R7081;
  wire [0:0] R7080;
  wire [0:0] R7079;
  wire [0:0] R7078;
  wire [0:0] R7077;
  wire [0:0] R7076;
  wire [0:0] R7075;
  wire [0:0] R7074;
  wire [0:0] R7073;
  wire [0:0] R7072;
  wire [0:0] R7071;
  wire [0:0] R7070;
  wire [0:0] R7069;
  wire [0:0] R7068;
  wire [0:0] R7067;
  wire [0:0] R7066;
  wire [0:0] R7065;
  wire [0:0] R7064;
  wire [0:0] R7063;
  wire [0:0] R7062;
  wire [0:0] R7061;
  wire [0:0] R7060;
  wire [0:0] R7059;
  wire [0:0] R7058;
  wire [0:0] R7057;
  wire [0:0] R7056;
  wire [0:0] R7055;
  wire [0:0] R7054;
  wire [0:0] R7053;
  wire [0:0] R7052;
  wire [0:0] R7051;
  wire [0:0] R7050;
  wire [0:0] R7049;
  wire [0:0] R7048;
  wire [0:0] R7047;
  wire [0:0] R7046;
  wire [0:0] R7045;
  wire [0:0] R7044;
  wire [0:0] R7043;
  wire [0:0] R7042;
  wire [0:0] R7041;
  wire [0:0] R7040;
  wire [0:0] R7039;
  wire [0:0] R7038;
  wire [0:0] R7037;
  wire [0:0] R7036;
  wire [0:0] R7035;
  wire [0:0] R7034;
  wire [0:0] R7033;
  wire [0:0] R7032;
  wire [0:0] R7031;
  wire [0:0] R7030;
  wire [0:0] R7029;
  wire [0:0] R7028;
  wire [63:0] R7027;
  wire [31:0] R7026;
  wire [31:0] R7025;
  wire [31:0] R7024;
  wire [31:0] R7023;
  wire [31:0] R7022;
  wire [31:0] R7021;
  wire [31:0] R7020;
  wire [31:0] R7019;
  wire [31:0] R7018;
  wire [31:0] R7017;
  wire [31:0] R7016;
  wire [31:0] R7015;
  wire [31:0] R7014;
  wire [31:0] R7013;
  wire [31:0] R7012;
  wire [31:0] R7011;
  wire [31:0] R7010;
  wire [31:0] R7009;
  wire [31:0] R7008;
  wire [31:0] R7007;
  wire [31:0] R7006;
  wire [31:0] R7005;
  wire [31:0] R7004;
  wire [31:0] R7003;
  wire [31:0] R7002;
  wire [31:0] R7001;
  wire [31:0] R7000;
  wire [31:0] R6999;
  wire [31:0] R6998;
  wire [31:0] R6997;
  wire [31:0] R6996;
  wire [31:0] R6995;
  wire [31:0] R6994;
  wire [31:0] R6993;
  wire [31:0] R6992;
  wire [31:0] R6991;
  wire [31:0] R6990;
  wire [31:0] R6989;
  wire [31:0] R6988;
  wire [31:0] R6987;
  wire [31:0] R6986;
  wire [31:0] R6985;
  wire [31:0] R6984;
  wire [31:0] R6983;
  wire [31:0] R6982;
  wire [31:0] R6981;
  wire [31:0] R6980;
  wire [31:0] R6979;
  wire [31:0] R6978;
  wire [31:0] R6977;
  wire [31:0] R6976;
  wire [31:0] R6975;
  wire [31:0] R6974;
  wire [31:0] R6973;
  wire [31:0] R6972;
  wire [31:0] R6971;
  wire [31:0] R6970;
  wire [31:0] R6969;
  wire [31:0] R6968;
  wire [31:0] R6967;
  wire [31:0] R6966;
  wire [31:0] R6965;
  wire [31:0] R6964;
  wire [31:0] R6963;
  wire [31:0] R6962;
  wire [31:0] R6961;
  wire [31:0] R6960;
  wire [31:0] R6959;
  wire [31:0] R6958;
  wire [31:0] R6957;
  wire [31:0] R6956;
  wire [31:0] R6955;
  wire [31:0] R6954;
  wire [31:0] R6953;
  wire [31:0] R6952;
  wire [31:0] R6951;
  wire [31:0] R6950;
  wire [31:0] R6949;
  wire [31:0] R6948;
  wire [31:0] R6947;
  wire [31:0] R6946;
  wire [31:0] R6945;
  wire [31:0] R6944;
  wire [31:0] R6943;
  wire [31:0] R6942;
  wire [31:0] R6941;
  wire [31:0] R6940;
  wire [31:0] R6939;
  wire [31:0] R6938;
  wire [63:0] R6937;
  wire [63:0] R6936;
  wire [63:0] R6935;
  wire [31:0] R6934;
  wire [31:0] R6933;
  wire [31:0] R6932;
  wire [31:0] R6931;
  wire [31:0] R6930;
  wire [31:0] R6929;
  wire [31:0] R6928;
  wire [31:0] R6927;
  wire [31:0] R6926;
  wire [31:0] R6925;
  wire [31:0] R6924;
  wire [31:0] R6923;
  wire [31:0] R6922;
  wire [31:0] R6921;
  wire [31:0] R6920;
  wire [31:0] R6919;
  wire [31:0] R6918;
  wire [31:0] R6917;
  wire [31:0] R6916;
  wire [31:0] R6915;
  wire [31:0] R6914;
  wire [31:0] R6913;
  wire [31:0] R6912;
  wire [31:0] R6911;
  wire [31:0] R6910;
  wire [31:0] R6909;
  wire [31:0] R6908;
  wire [31:0] R6907;
  wire [31:0] R6906;
  wire [31:0] R6905;
  wire [31:0] R6904;
  wire [31:0] R6903;
  wire [31:0] R6902;
  wire [31:0] R6901;
  wire [31:0] R6900;
  wire [31:0] R6899;
  wire [31:0] R6898;
  wire [31:0] R6897;
  wire [31:0] R6896;
  wire [31:0] R6895;
  wire [31:0] R6894;
  wire [31:0] R6893;
  wire [31:0] R6892;
  wire [31:0] R6891;
  wire [31:0] R6890;
  wire [31:0] R6889;
  wire [31:0] R6888;
  wire [31:0] R6887;
  wire [31:0] R6886;
  wire [31:0] R6885;
  wire [31:0] R6884;
  wire [31:0] R6883;
  wire [31:0] R6882;
  wire [31:0] R6881;
  wire [31:0] R6880;
  wire [31:0] R6879;
  wire [31:0] R6878;
  wire [31:0] R6877;
  wire [31:0] R6876;
  wire [31:0] R6875;
  wire [31:0] R6874;
  wire [31:0] R6873;
  wire [31:0] R6872;
  wire [31:0] R6871;
  wire [31:0] R6870;
  wire [31:0] R6869;
  wire [31:0] R6868;
  wire [31:0] R6867;
  wire [31:0] R6866;
  wire [31:0] R6865;
  wire [31:0] R6864;
  wire [31:0] R6863;
  wire [31:0] R6862;
  wire [31:0] R6861;
  wire [31:0] R6860;
  wire [31:0] R6859;
  wire [31:0] R6858;
  wire [31:0] R6857;
  wire [31:0] R6856;
  wire [31:0] R6855;
  wire [31:0] R6854;
  wire [31:0] R6853;
  wire [31:0] R6852;
  wire [31:0] R6851;
  wire [31:0] R6850;
  wire [31:0] R6849;
  wire [31:0] R6848;
  wire [31:0] R6847;
  wire [31:0] R6846;
  wire [31:0] R6845;
  wire [31:0] R6844;
  wire [31:0] R6843;
  wire [31:0] R6842;
  wire [31:0] R6841;
  wire [31:0] R6840;
  wire [31:0] R6839;
  wire [63:0] R6838;
  wire [31:0] R6837;
  wire [31:0] R6836;
  wire [63:0] R6835;
  wire [31:0] R6834;
  wire [63:0] R6833;
  wire [63:0] R6832;
  wire [63:0] R6831;
  wire [63:0] R6830;
  wire [63:0] R6829;
  wire [63:0] R6828;
  wire [31:0] R6827;
  wire [63:0] R6826;
  wire [63:0] R6825;
  wire [63:0] R6824;
  wire [63:0] R6823;
  wire [63:0] R6822;
  wire [63:0] R6821;
  wire [63:0] R6820;
  wire [31:0] R6819;
  wire [31:0] R6818;
  wire [31:0] R6817;
  wire [63:0] R6816;
  wire [63:0] R6815;
  wire [63:0] R6814;
  wire [63:0] R6813;
  wire [63:0] R6812;
  wire [63:0] R6811;
  wire [63:0] R6810;
  wire [63:0] R6809;
  wire [63:0] R6808;
  wire [63:0] R6807;
  wire [63:0] R6806;
  wire [63:0] R6805;
  wire [63:0] R6804;
  wire [63:0] R6803;
  wire [63:0] R6802;
  wire [63:0] R6801;
  wire [63:0] R6800;
  wire [63:0] R6799;
  wire [63:0] R6798;
  wire [63:0] R6797;
  wire [63:0] R6796;
  wire [63:0] R6795;
  wire [63:0] R6794;
  wire [63:0] R6793;
  wire [0:0] R6792;
  wire [0:0] R6791;
  wire [0:0] R6790;
  wire [0:0] R6789;
  wire [0:0] R6788;
  wire [0:0] R6787;
  wire [0:0] R6786;
  wire [0:0] R6785;
  wire [0:0] R6784;
  wire [0:0] R6783;
  wire [0:0] R6782;
  wire [0:0] R6781;
  wire [0:0] R6780;
  wire [0:0] R6779;
  wire [0:0] R6778;
  wire [0:0] R6777;
  wire [0:0] R6776;
  wire [0:0] R6775;
  wire [0:0] R6774;
  wire [0:0] R6773;
  wire [0:0] R6772;
  wire [0:0] R6771;
  wire [0:0] R6770;
  wire [0:0] R6769;
  wire [0:0] R6768;
  wire [0:0] R6767;
  wire [0:0] R6766;
  wire [0:0] R6765;
  wire [0:0] R6764;
  wire [0:0] R6763;
  wire [0:0] R6762;
  wire [0:0] R6761;
  wire [0:0] R6760;
  wire [0:0] R6759;
  wire [0:0] R6758;
  wire [0:0] R6757;
  wire [0:0] R6756;
  wire [0:0] R6755;
  wire [0:0] R6754;
  wire [0:0] R6753;
  wire [0:0] R6752;
  wire [0:0] R6751;
  wire [0:0] R6750;
  wire [0:0] R6749;
  wire [0:0] R6748;
  wire [0:0] R6747;
  wire [0:0] R6746;
  wire [0:0] R6745;
  wire [0:0] R6744;
  wire [0:0] R6743;
  wire [0:0] R6742;
  wire [0:0] R6741;
  wire [0:0] R6740;
  wire [0:0] R6739;
  wire [0:0] R6738;
  wire [0:0] R6737;
  wire [0:0] R6736;
  wire [0:0] R6735;
  wire [0:0] R6734;
  wire [0:0] R6733;
  wire [0:0] R6732;
  wire [0:0] R6731;
  wire [0:0] R6730;
  wire [0:0] R6729;
  wire [0:0] R6728;
  wire [0:0] R6727;
  wire [0:0] R6726;
  wire [0:0] R6725;
  wire [0:0] R6724;
  wire [0:0] R6723;
  wire [0:0] R6722;
  wire [0:0] R6721;
  wire [0:0] R6720;
  wire [0:0] R6719;
  wire [0:0] R6718;
  wire [0:0] R6717;
  wire [0:0] R6716;
  wire [0:0] R6715;
  wire [0:0] R6714;
  wire [0:0] R6713;
  wire [0:0] R6712;
  wire [0:0] R6711;
  wire [0:0] R6710;
  wire [0:0] R6709;
  wire [0:0] R6708;
  wire [0:0] R6707;
  wire [0:0] R6706;
  wire [0:0] R6705;
  wire [0:0] R6704;
  wire [0:0] R6703;
  wire [0:0] R6702;
  wire [0:0] R6701;
  wire [0:0] R6700;
  wire [0:0] R6699;
  wire [0:0] R6698;
  wire [0:0] R6697;
  wire [0:0] R6696;
  wire [0:0] R6695;
  wire [0:0] R6694;
  wire [0:0] R6693;
  wire [0:0] R6692;
  wire [0:0] R6691;
  wire [0:0] R6690;
  wire [0:0] R6689;
  wire [0:0] R6688;
  wire [0:0] R6687;
  wire [0:0] R6686;
  wire [0:0] R6685;
  wire [0:0] R6684;
  wire [63:0] R6683;
  wire [31:0] R6682;
  wire [31:0] R6681;
  wire [31:0] R6680;
  wire [31:0] R6679;
  wire [31:0] R6678;
  wire [31:0] R6677;
  wire [31:0] R6676;
  wire [31:0] R6675;
  wire [31:0] R6674;
  wire [31:0] R6673;
  wire [31:0] R6672;
  wire [31:0] R6671;
  wire [31:0] R6670;
  wire [31:0] R6669;
  wire [31:0] R6668;
  wire [31:0] R6667;
  wire [31:0] R6666;
  wire [31:0] R6665;
  wire [31:0] R6664;
  wire [31:0] R6663;
  wire [31:0] R6662;
  wire [31:0] R6661;
  wire [31:0] R6660;
  wire [31:0] R6659;
  wire [31:0] R6658;
  wire [31:0] R6657;
  wire [31:0] R6656;
  wire [31:0] R6655;
  wire [31:0] R6654;
  wire [31:0] R6653;
  wire [31:0] R6652;
  wire [31:0] R6651;
  wire [31:0] R6650;
  wire [31:0] R6649;
  wire [31:0] R6648;
  wire [31:0] R6647;
  wire [31:0] R6646;
  wire [31:0] R6645;
  wire [31:0] R6644;
  wire [31:0] R6643;
  wire [31:0] R6642;
  wire [31:0] R6641;
  wire [31:0] R6640;
  wire [31:0] R6639;
  wire [31:0] R6638;
  wire [31:0] R6637;
  wire [31:0] R6636;
  wire [31:0] R6635;
  wire [31:0] R6634;
  wire [31:0] R6633;
  wire [31:0] R6632;
  wire [31:0] R6631;
  wire [31:0] R6630;
  wire [31:0] R6629;
  wire [31:0] R6628;
  wire [31:0] R6627;
  wire [31:0] R6626;
  wire [31:0] R6625;
  wire [31:0] R6624;
  wire [31:0] R6623;
  wire [31:0] R6622;
  wire [31:0] R6621;
  wire [31:0] R6620;
  wire [31:0] R6619;
  wire [31:0] R6618;
  wire [31:0] R6617;
  wire [31:0] R6616;
  wire [31:0] R6615;
  wire [31:0] R6614;
  wire [31:0] R6613;
  wire [31:0] R6612;
  wire [31:0] R6611;
  wire [31:0] R6610;
  wire [31:0] R6609;
  wire [31:0] R6608;
  wire [31:0] R6607;
  wire [31:0] R6606;
  wire [31:0] R6605;
  wire [31:0] R6604;
  wire [31:0] R6603;
  wire [31:0] R6602;
  wire [31:0] R6601;
  wire [31:0] R6600;
  wire [31:0] R6599;
  wire [31:0] R6598;
  wire [31:0] R6597;
  wire [31:0] R6596;
  wire [31:0] R6595;
  wire [31:0] R6594;
  wire [31:0] R6593;
  wire [31:0] R6592;
  wire [31:0] R6591;
  wire [31:0] R6590;
  wire [31:0] R6589;
  wire [31:0] R6588;
  wire [31:0] R6587;
  wire [31:0] R6586;
  wire [31:0] R6585;
  wire [31:0] R6584;
  wire [31:0] R6583;
  wire [31:0] R6582;
  wire [31:0] R6581;
  wire [31:0] R6580;
  wire [63:0] R6579;
  wire [63:0] R6578;
  wire [63:0] R6577;
  wire [31:0] R6576;
  wire [31:0] R6575;
  wire [31:0] R6574;
  wire [31:0] R6573;
  wire [31:0] R6572;
  wire [31:0] R6571;
  wire [31:0] R6570;
  wire [31:0] R6569;
  wire [31:0] R6568;
  wire [31:0] R6567;
  wire [31:0] R6566;
  wire [31:0] R6565;
  wire [31:0] R6564;
  wire [31:0] R6563;
  wire [31:0] R6562;
  wire [31:0] R6561;
  wire [31:0] R6560;
  wire [31:0] R6559;
  wire [31:0] R6558;
  wire [31:0] R6557;
  wire [31:0] R6556;
  wire [31:0] R6555;
  wire [31:0] R6554;
  wire [31:0] R6553;
  wire [31:0] R6552;
  wire [31:0] R6551;
  wire [31:0] R6550;
  wire [31:0] R6549;
  wire [31:0] R6548;
  wire [31:0] R6547;
  wire [31:0] R6546;
  wire [31:0] R6545;
  wire [31:0] R6544;
  wire [31:0] R6543;
  wire [31:0] R6542;
  wire [31:0] R6541;
  wire [31:0] R6540;
  wire [31:0] R6539;
  wire [31:0] R6538;
  wire [31:0] R6537;
  wire [31:0] R6536;
  wire [31:0] R6535;
  wire [31:0] R6534;
  wire [31:0] R6533;
  wire [31:0] R6532;
  wire [31:0] R6531;
  wire [31:0] R6530;
  wire [31:0] R6529;
  wire [31:0] R6528;
  wire [31:0] R6527;
  wire [31:0] R6526;
  wire [31:0] R6525;
  wire [31:0] R6524;
  wire [31:0] R6523;
  wire [31:0] R6522;
  wire [31:0] R6521;
  wire [31:0] R6520;
  wire [31:0] R6519;
  wire [31:0] R6518;
  wire [31:0] R6517;
  wire [31:0] R6516;
  wire [31:0] R6515;
  wire [31:0] R6514;
  wire [31:0] R6513;
  wire [31:0] R6512;
  wire [31:0] R6511;
  wire [31:0] R6510;
  wire [31:0] R6509;
  wire [31:0] R6508;
  wire [31:0] R6507;
  wire [31:0] R6506;
  wire [31:0] R6505;
  wire [31:0] R6504;
  wire [31:0] R6503;
  wire [31:0] R6502;
  wire [31:0] R6501;
  wire [31:0] R6500;
  wire [31:0] R6499;
  wire [31:0] R6498;
  wire [31:0] R6497;
  wire [31:0] R6496;
  wire [31:0] R6495;
  wire [31:0] R6494;
  wire [31:0] R6493;
  wire [31:0] R6492;
  wire [31:0] R6491;
  wire [31:0] R6490;
  wire [31:0] R6489;
  wire [31:0] R6488;
  wire [31:0] R6487;
  wire [31:0] R6486;
  wire [31:0] R6485;
  wire [31:0] R6484;
  wire [31:0] R6483;
  wire [31:0] R6482;
  wire [31:0] R6481;
  wire [31:0] R6480;
  wire [31:0] R6479;
  wire [31:0] R6478;
  wire [31:0] R6477;
  wire [31:0] R6476;
  wire [31:0] R6475;
  wire [31:0] R6474;
  wire [31:0] R6473;
  wire [31:0] R6472;
  wire [31:0] R6471;
  wire [31:0] R6470;
  wire [31:0] R6469;
  wire [31:0] R6468;
  wire [31:0] R6467;
  wire [63:0] R6466;
  wire [31:0] R6465;
  wire [31:0] R6464;
  wire [63:0] R6463;
  wire [31:0] R6462;
  wire [63:0] R6461;
  wire [63:0] R6460;
  wire [63:0] R6459;
  wire [63:0] R6458;
  wire [63:0] R6457;
  wire [63:0] R6456;
  wire [31:0] R6455;
  wire [63:0] R6454;
  wire [63:0] R6453;
  wire [63:0] R6452;
  wire [63:0] R6451;
  wire [63:0] R6450;
  wire [63:0] R6449;
  wire [63:0] R6448;
  wire [31:0] R6447;
  wire [31:0] R6446;
  wire [31:0] R6445;
  wire [63:0] R6444;
  wire [63:0] R6443;
  wire [63:0] R6442;
  wire [63:0] R6441;
  wire [63:0] R6440;
  wire [63:0] R6439;
  wire [63:0] R6438;
  wire [63:0] R6437;
  wire [63:0] R6436;
  wire [63:0] R6435;
  wire [63:0] R6434;
  wire [63:0] R6433;
  wire [63:0] R6432;
  wire [63:0] R6431;
  wire [63:0] R6430;
  wire [63:0] R6429;
  wire [63:0] R6428;
  wire [63:0] R6427;
  wire [63:0] R6426;
  wire [63:0] R6425;
  wire [63:0] R6424;
  wire [63:0] R6423;
  wire [63:0] R6422;
  wire [63:0] R6421;
  wire [0:0] R6420;
  wire [0:0] R6419;
  wire [0:0] R6418;
  wire [0:0] R6417;
  wire [0:0] R6416;
  wire [0:0] R6415;
  wire [0:0] R6414;
  wire [0:0] R6413;
  wire [0:0] R6412;
  wire [0:0] R6411;
  wire [0:0] R6410;
  wire [0:0] R6409;
  wire [0:0] R6408;
  wire [0:0] R6407;
  wire [0:0] R6406;
  wire [0:0] R6405;
  wire [0:0] R6404;
  wire [0:0] R6403;
  wire [0:0] R6402;
  wire [0:0] R6401;
  wire [0:0] R6400;
  wire [0:0] R6399;
  wire [0:0] R6398;
  wire [0:0] R6397;
  wire [0:0] R6396;
  wire [0:0] R6395;
  wire [0:0] R6394;
  wire [0:0] R6393;
  wire [0:0] R6392;
  wire [0:0] R6391;
  wire [0:0] R6390;
  wire [0:0] R6389;
  wire [0:0] R6388;
  wire [0:0] R6387;
  wire [0:0] R6386;
  wire [0:0] R6385;
  wire [0:0] R6384;
  wire [0:0] R6383;
  wire [0:0] R6382;
  wire [0:0] R6381;
  wire [0:0] R6380;
  wire [0:0] R6379;
  wire [0:0] R6378;
  wire [0:0] R6377;
  wire [0:0] R6376;
  wire [0:0] R6375;
  wire [0:0] R6374;
  wire [0:0] R6373;
  wire [0:0] R6372;
  wire [0:0] R6371;
  wire [0:0] R6370;
  wire [0:0] R6369;
  wire [0:0] R6368;
  wire [0:0] R6367;
  wire [0:0] R6366;
  wire [0:0] R6365;
  wire [0:0] R6364;
  wire [0:0] R6363;
  wire [0:0] R6362;
  wire [0:0] R6361;
  wire [0:0] R6360;
  wire [0:0] R6359;
  wire [0:0] R6358;
  wire [0:0] R6357;
  wire [0:0] R6356;
  wire [0:0] R6355;
  wire [0:0] R6354;
  wire [0:0] R6353;
  wire [0:0] R6352;
  wire [0:0] R6351;
  wire [0:0] R6350;
  wire [0:0] R6349;
  wire [0:0] R6348;
  wire [0:0] R6347;
  wire [0:0] R6346;
  wire [0:0] R6345;
  wire [0:0] R6344;
  wire [0:0] R6343;
  wire [0:0] R6342;
  wire [0:0] R6341;
  wire [0:0] R6340;
  wire [0:0] R6339;
  wire [0:0] R6338;
  wire [0:0] R6337;
  wire [0:0] R6336;
  wire [0:0] R6335;
  wire [0:0] R6334;
  wire [0:0] R6333;
  wire [0:0] R6332;
  wire [0:0] R6331;
  wire [0:0] R6330;
  wire [0:0] R6329;
  wire [0:0] R6328;
  wire [0:0] R6327;
  wire [0:0] R6326;
  wire [0:0] R6325;
  wire [0:0] R6324;
  wire [0:0] R6323;
  wire [0:0] R6322;
  wire [0:0] R6321;
  wire [0:0] R6320;
  wire [0:0] R6319;
  wire [0:0] R6318;
  wire [0:0] R6317;
  wire [0:0] R6316;
  wire [0:0] R6315;
  wire [0:0] R6314;
  wire [0:0] R6313;
  wire [0:0] R6312;
  wire [0:0] R6311;
  wire [0:0] R6310;
  wire [0:0] R6309;
  wire [0:0] R6308;
  wire [0:0] R6307;
  wire [0:0] R6306;
  wire [0:0] R6305;
  wire [0:0] R6304;
  wire [0:0] R6303;
  wire [0:0] R6302;
  wire [0:0] R6301;
  wire [0:0] R6300;
  wire [0:0] R6299;
  wire [0:0] R6298;
  wire [0:0] R6297;
  wire [63:0] R6296;
  wire [31:0] R6295;
  wire [31:0] R6294;
  wire [31:0] R6293;
  wire [31:0] R6292;
  wire [31:0] R6291;
  wire [31:0] R6290;
  wire [31:0] R6289;
  wire [31:0] R6288;
  wire [31:0] R6287;
  wire [31:0] R6286;
  wire [31:0] R6285;
  wire [31:0] R6284;
  wire [31:0] R6283;
  wire [31:0] R6282;
  wire [31:0] R6281;
  wire [31:0] R6280;
  wire [31:0] R6279;
  wire [31:0] R6278;
  wire [31:0] R6277;
  wire [31:0] R6276;
  wire [31:0] R6275;
  wire [31:0] R6274;
  wire [31:0] R6273;
  wire [31:0] R6272;
  wire [31:0] R6271;
  wire [31:0] R6270;
  wire [31:0] R6269;
  wire [31:0] R6268;
  wire [31:0] R6267;
  wire [31:0] R6266;
  wire [31:0] R6265;
  wire [31:0] R6264;
  wire [31:0] R6263;
  wire [31:0] R6262;
  wire [31:0] R6261;
  wire [31:0] R6260;
  wire [31:0] R6259;
  wire [31:0] R6258;
  wire [31:0] R6257;
  wire [31:0] R6256;
  wire [31:0] R6255;
  wire [31:0] R6254;
  wire [31:0] R6253;
  wire [31:0] R6252;
  wire [31:0] R6251;
  wire [31:0] R6250;
  wire [31:0] R6249;
  wire [31:0] R6248;
  wire [31:0] R6247;
  wire [31:0] R6246;
  wire [31:0] R6245;
  wire [31:0] R6244;
  wire [31:0] R6243;
  wire [31:0] R6242;
  wire [31:0] R6241;
  wire [31:0] R6240;
  wire [31:0] R6239;
  wire [31:0] R6238;
  wire [31:0] R6237;
  wire [31:0] R6236;
  wire [31:0] R6235;
  wire [31:0] R6234;
  wire [31:0] R6233;
  wire [31:0] R6232;
  wire [31:0] R6231;
  wire [31:0] R6230;
  wire [31:0] R6229;
  wire [31:0] R6228;
  wire [31:0] R6227;
  wire [31:0] R6226;
  wire [31:0] R6225;
  wire [31:0] R6224;
  wire [31:0] R6223;
  wire [31:0] R6222;
  wire [31:0] R6221;
  wire [31:0] R6220;
  wire [31:0] R6219;
  wire [31:0] R6218;
  wire [31:0] R6217;
  wire [31:0] R6216;
  wire [31:0] R6215;
  wire [31:0] R6214;
  wire [31:0] R6213;
  wire [31:0] R6212;
  wire [31:0] R6211;
  wire [31:0] R6210;
  wire [31:0] R6209;
  wire [31:0] R6208;
  wire [31:0] R6207;
  wire [31:0] R6206;
  wire [31:0] R6205;
  wire [31:0] R6204;
  wire [31:0] R6203;
  wire [31:0] R6202;
  wire [31:0] R6201;
  wire [31:0] R6200;
  wire [31:0] R6199;
  wire [31:0] R6198;
  wire [31:0] R6197;
  wire [31:0] R6196;
  wire [31:0] R6195;
  wire [31:0] R6194;
  wire [31:0] R6193;
  wire [31:0] R6192;
  wire [31:0] R6191;
  wire [31:0] R6190;
  wire [31:0] R6189;
  wire [31:0] R6188;
  wire [31:0] R6187;
  wire [31:0] R6186;
  wire [31:0] R6185;
  wire [31:0] R6184;
  wire [31:0] R6183;
  wire [31:0] R6182;
  wire [31:0] R6181;
  wire [31:0] R6180;
  wire [31:0] R6179;
  wire [63:0] R6178;
  wire [63:0] R6177;
  wire [63:0] R6176;
  wire [31:0] R6175;
  wire [31:0] R6174;
  wire [31:0] R6173;
  wire [31:0] R6172;
  wire [31:0] R6171;
  wire [31:0] R6170;
  wire [31:0] R6169;
  wire [31:0] R6168;
  wire [31:0] R6167;
  wire [31:0] R6166;
  wire [31:0] R6165;
  wire [31:0] R6164;
  wire [31:0] R6163;
  wire [31:0] R6162;
  wire [31:0] R6161;
  wire [31:0] R6160;
  wire [31:0] R6159;
  wire [31:0] R6158;
  wire [31:0] R6157;
  wire [31:0] R6156;
  wire [31:0] R6155;
  wire [31:0] R6154;
  wire [31:0] R6153;
  wire [31:0] R6152;
  wire [31:0] R6151;
  wire [31:0] R6150;
  wire [31:0] R6149;
  wire [31:0] R6148;
  wire [31:0] R6147;
  wire [31:0] R6146;
  wire [31:0] R6145;
  wire [31:0] R6144;
  wire [31:0] R6143;
  wire [31:0] R6142;
  wire [31:0] R6141;
  wire [31:0] R6140;
  wire [31:0] R6139;
  wire [31:0] R6138;
  wire [31:0] R6137;
  wire [31:0] R6136;
  wire [31:0] R6135;
  wire [31:0] R6134;
  wire [31:0] R6133;
  wire [31:0] R6132;
  wire [31:0] R6131;
  wire [31:0] R6130;
  wire [31:0] R6129;
  wire [31:0] R6128;
  wire [31:0] R6127;
  wire [31:0] R6126;
  wire [31:0] R6125;
  wire [31:0] R6124;
  wire [31:0] R6123;
  wire [31:0] R6122;
  wire [31:0] R6121;
  wire [31:0] R6120;
  wire [31:0] R6119;
  wire [31:0] R6118;
  wire [31:0] R6117;
  wire [31:0] R6116;
  wire [31:0] R6115;
  wire [31:0] R6114;
  wire [31:0] R6113;
  wire [31:0] R6112;
  wire [31:0] R6111;
  wire [31:0] R6110;
  wire [31:0] R6109;
  wire [31:0] R6108;
  wire [31:0] R6107;
  wire [31:0] R6106;
  wire [31:0] R6105;
  wire [31:0] R6104;
  wire [31:0] R6103;
  wire [31:0] R6102;
  wire [31:0] R6101;
  wire [31:0] R6100;
  wire [31:0] R6099;
  wire [31:0] R6098;
  wire [31:0] R6097;
  wire [31:0] R6096;
  wire [31:0] R6095;
  wire [31:0] R6094;
  wire [31:0] R6093;
  wire [31:0] R6092;
  wire [31:0] R6091;
  wire [31:0] R6090;
  wire [31:0] R6089;
  wire [31:0] R6088;
  wire [31:0] R6087;
  wire [31:0] R6086;
  wire [31:0] R6085;
  wire [31:0] R6084;
  wire [31:0] R6083;
  wire [31:0] R6082;
  wire [31:0] R6081;
  wire [31:0] R6080;
  wire [31:0] R6079;
  wire [31:0] R6078;
  wire [31:0] R6077;
  wire [31:0] R6076;
  wire [31:0] R6075;
  wire [31:0] R6074;
  wire [31:0] R6073;
  wire [31:0] R6072;
  wire [31:0] R6071;
  wire [31:0] R6070;
  wire [31:0] R6069;
  wire [31:0] R6068;
  wire [31:0] R6067;
  wire [31:0] R6066;
  wire [31:0] R6065;
  wire [31:0] R6064;
  wire [31:0] R6063;
  wire [31:0] R6062;
  wire [31:0] R6061;
  wire [31:0] R6060;
  wire [31:0] R6059;
  wire [31:0] R6058;
  wire [31:0] R6057;
  wire [31:0] R6056;
  wire [31:0] R6055;
  wire [31:0] R6054;
  wire [31:0] R6053;
  wire [31:0] R6052;
  wire [31:0] R6051;
  wire [31:0] R6050;
  wire [63:0] R6049;
  wire [31:0] R6048;
  wire [63:0] R6047;
  wire [63:0] R6046;
  wire [63:0] R6045;
  wire [63:0] R6044;
  wire [63:0] R6043;
  wire [63:0] R6042;
  wire [31:0] R6041;
  wire [63:0] R6040;
  wire [63:0] R6039;
  wire [63:0] R6038;
  wire [63:0] R6037;
  wire [63:0] R6036;
  wire [63:0] R6035;
  wire [63:0] R6034;
  wire [31:0] R6033;
  wire [31:0] R6032;
  wire [31:0] R6031;
  wire [63:0] R6030;
  wire [63:0] R6029;
  wire [63:0] R6028;
  wire [63:0] R6027;
  wire [63:0] R6026;
  wire [63:0] R6025;
  wire [63:0] R6024;
  wire [63:0] R6023;
  wire [63:0] R6022;
  wire [63:0] R6021;
  wire [63:0] R6020;
  wire [63:0] R6019;
  wire [63:0] R6018;
  wire [63:0] R6017;
  wire [63:0] R6016;
  wire [63:0] R6015;
  wire [63:0] R6014;
  wire [63:0] R6013;
  wire [63:0] R6012;
  wire [63:0] R6011;
  wire [63:0] R6010;
  wire [63:0] R6009;
  wire [63:0] R6008;
  wire [63:0] R6007;
  wire [0:0] R6006;
  wire [0:0] R6005;
  wire [0:0] R6004;
  wire [0:0] R6003;
  wire [0:0] R6002;
  wire [0:0] R6001;
  wire [0:0] R6000;
  wire [0:0] R5999;
  wire [0:0] R5998;
  wire [0:0] R5997;
  wire [0:0] R5996;
  wire [0:0] R5995;
  wire [0:0] R5994;
  wire [0:0] R5993;
  wire [0:0] R5992;
  wire [0:0] R5991;
  wire [0:0] R5990;
  wire [0:0] R5989;
  wire [0:0] R5988;
  wire [0:0] R5987;
  wire [0:0] R5986;
  wire [0:0] R5985;
  wire [0:0] R5984;
  wire [0:0] R5983;
  wire [0:0] R5982;
  wire [0:0] R5981;
  wire [0:0] R5980;
  wire [0:0] R5979;
  wire [0:0] R5978;
  wire [0:0] R5977;
  wire [0:0] R5976;
  wire [0:0] R5975;
  wire [0:0] R5974;
  wire [0:0] R5973;
  wire [0:0] R5972;
  wire [0:0] R5971;
  wire [0:0] R5970;
  wire [0:0] R5969;
  wire [0:0] R5968;
  wire [0:0] R5967;
  wire [0:0] R5966;
  wire [0:0] R5965;
  wire [0:0] R5964;
  wire [0:0] R5963;
  wire [0:0] R5962;
  wire [0:0] R5961;
  wire [0:0] R5960;
  wire [0:0] R5959;
  wire [0:0] R5958;
  wire [0:0] R5957;
  wire [0:0] R5956;
  wire [0:0] R5955;
  wire [0:0] R5954;
  wire [0:0] R5953;
  wire [0:0] R5952;
  wire [0:0] R5951;
  wire [0:0] R5950;
  wire [0:0] R5949;
  wire [0:0] R5948;
  wire [0:0] R5947;
  wire [0:0] R5946;
  wire [0:0] R5945;
  wire [0:0] R5944;
  wire [0:0] R5943;
  wire [0:0] R5942;
  wire [0:0] R5941;
  wire [0:0] R5940;
  wire [0:0] R5939;
  wire [0:0] R5938;
  wire [0:0] R5937;
  wire [0:0] R5936;
  wire [0:0] R5935;
  wire [0:0] R5934;
  wire [0:0] R5933;
  wire [0:0] R5932;
  wire [0:0] R5931;
  wire [0:0] R5930;
  wire [0:0] R5929;
  wire [0:0] R5928;
  wire [0:0] R5927;
  wire [0:0] R5926;
  wire [0:0] R5925;
  wire [0:0] R5924;
  wire [0:0] R5923;
  wire [0:0] R5922;
  wire [0:0] R5921;
  wire [0:0] R5920;
  wire [0:0] R5919;
  wire [0:0] R5918;
  wire [0:0] R5917;
  wire [0:0] R5916;
  wire [0:0] R5915;
  wire [0:0] R5914;
  wire [0:0] R5913;
  wire [0:0] R5912;
  wire [0:0] R5911;
  wire [0:0] R5910;
  wire [0:0] R5909;
  wire [0:0] R5908;
  wire [0:0] R5907;
  wire [0:0] R5906;
  wire [0:0] R5905;
  wire [0:0] R5904;
  wire [0:0] R5903;
  wire [0:0] R5902;
  wire [0:0] R5901;
  wire [0:0] R5900;
  wire [0:0] R5899;
  wire [0:0] R5898;
  wire [0:0] R5897;
  wire [0:0] R5896;
  wire [0:0] R5895;
  wire [0:0] R5894;
  wire [0:0] R5893;
  wire [0:0] R5892;
  wire [0:0] R5891;
  wire [0:0] R5890;
  wire [0:0] R5889;
  wire [0:0] R5888;
  wire [0:0] R5887;
  wire [0:0] R5886;
  wire [0:0] R5885;
  wire [0:0] R5884;
  wire [0:0] R5883;
  wire [0:0] R5882;
  wire [0:0] R5881;
  wire [0:0] R5880;
  wire [0:0] R5879;
  wire [0:0] R5878;
  wire [0:0] R5877;
  wire [0:0] R5876;
  wire [0:0] R5875;
  wire [0:0] R5874;
  wire [0:0] R5873;
  wire [0:0] R5872;
  wire [0:0] R5871;
  wire [0:0] R5870;
  wire [0:0] R5869;
  wire [63:0] R5868;
  wire [31:0] R5867;
  wire [31:0] R5866;
  wire [31:0] R5865;
  wire [31:0] R5864;
  wire [31:0] R5863;
  wire [31:0] R5862;
  wire [31:0] R5861;
  wire [31:0] R5860;
  wire [31:0] R5859;
  wire [31:0] R5858;
  wire [31:0] R5857;
  wire [31:0] R5856;
  wire [31:0] R5855;
  wire [31:0] R5854;
  wire [31:0] R5853;
  wire [31:0] R5852;
  wire [31:0] R5851;
  wire [31:0] R5850;
  wire [31:0] R5849;
  wire [31:0] R5848;
  wire [31:0] R5847;
  wire [31:0] R5846;
  wire [31:0] R5845;
  wire [31:0] R5844;
  wire [31:0] R5843;
  wire [31:0] R5842;
  wire [31:0] R5841;
  wire [31:0] R5840;
  wire [31:0] R5839;
  wire [31:0] R5838;
  wire [31:0] R5837;
  wire [31:0] R5836;
  wire [31:0] R5835;
  wire [31:0] R5834;
  wire [31:0] R5833;
  wire [31:0] R5832;
  wire [31:0] R5831;
  wire [31:0] R5830;
  wire [31:0] R5829;
  wire [31:0] R5828;
  wire [31:0] R5827;
  wire [31:0] R5826;
  wire [31:0] R5825;
  wire [31:0] R5824;
  wire [31:0] R5823;
  wire [31:0] R5822;
  wire [31:0] R5821;
  wire [31:0] R5820;
  wire [31:0] R5819;
  wire [31:0] R5818;
  wire [31:0] R5817;
  wire [31:0] R5816;
  wire [31:0] R5815;
  wire [31:0] R5814;
  wire [31:0] R5813;
  wire [31:0] R5812;
  wire [31:0] R5811;
  wire [31:0] R5810;
  wire [31:0] R5809;
  wire [31:0] R5808;
  wire [31:0] R5807;
  wire [31:0] R5806;
  wire [31:0] R5805;
  wire [31:0] R5804;
  wire [31:0] R5803;
  wire [31:0] R5802;
  wire [31:0] R5801;
  wire [31:0] R5800;
  wire [31:0] R5799;
  wire [31:0] R5798;
  wire [31:0] R5797;
  wire [31:0] R5796;
  wire [31:0] R5795;
  wire [31:0] R5794;
  wire [31:0] R5793;
  wire [31:0] R5792;
  wire [31:0] R5791;
  wire [31:0] R5790;
  wire [31:0] R5789;
  wire [31:0] R5788;
  wire [31:0] R5787;
  wire [31:0] R5786;
  wire [31:0] R5785;
  wire [31:0] R5784;
  wire [31:0] R5783;
  wire [31:0] R5782;
  wire [31:0] R5781;
  wire [31:0] R5780;
  wire [31:0] R5779;
  wire [31:0] R5778;
  wire [31:0] R5777;
  wire [31:0] R5776;
  wire [31:0] R5775;
  wire [31:0] R5774;
  wire [31:0] R5773;
  wire [31:0] R5772;
  wire [31:0] R5771;
  wire [31:0] R5770;
  wire [31:0] R5769;
  wire [31:0] R5768;
  wire [31:0] R5767;
  wire [31:0] R5766;
  wire [31:0] R5765;
  wire [31:0] R5764;
  wire [31:0] R5763;
  wire [31:0] R5762;
  wire [31:0] R5761;
  wire [31:0] R5760;
  wire [31:0] R5759;
  wire [31:0] R5758;
  wire [31:0] R5757;
  wire [31:0] R5756;
  wire [31:0] R5755;
  wire [31:0] R5754;
  wire [31:0] R5753;
  wire [31:0] R5752;
  wire [31:0] R5751;
  wire [31:0] R5750;
  wire [31:0] R5749;
  wire [31:0] R5748;
  wire [31:0] R5747;
  wire [31:0] R5746;
  wire [31:0] R5745;
  wire [31:0] R5744;
  wire [31:0] R5743;
  wire [31:0] R5742;
  wire [31:0] R5741;
  wire [31:0] R5740;
  wire [31:0] R5739;
  wire [31:0] R5738;
  wire [31:0] R5737;
  wire [31:0] R5736;
  wire [63:0] R5735;
  wire [63:0] R5734;
  wire [63:0] R5733;
  wire [31:0] R5732;
  wire [31:0] R5731;
  wire [31:0] R5730;
  wire [31:0] R5729;
  wire [31:0] R5728;
  wire [31:0] R5727;
  wire [31:0] R5726;
  wire [31:0] R5725;
  wire [31:0] R5724;
  wire [31:0] R5723;
  wire [31:0] R5722;
  wire [31:0] R5721;
  wire [31:0] R5720;
  wire [31:0] R5719;
  wire [31:0] R5718;
  wire [31:0] R5717;
  wire [31:0] R5716;
  wire [31:0] R5715;
  wire [31:0] R5714;
  wire [31:0] R5713;
  wire [31:0] R5712;
  wire [31:0] R5711;
  wire [31:0] R5710;
  wire [31:0] R5709;
  wire [31:0] R5708;
  wire [31:0] R5707;
  wire [31:0] R5706;
  wire [31:0] R5705;
  wire [31:0] R5704;
  wire [31:0] R5703;
  wire [31:0] R5702;
  wire [31:0] R5701;
  wire [31:0] R5700;
  wire [31:0] R5699;
  wire [31:0] R5698;
  wire [31:0] R5697;
  wire [31:0] R5696;
  wire [31:0] R5695;
  wire [31:0] R5694;
  wire [31:0] R5693;
  wire [31:0] R5692;
  wire [31:0] R5691;
  wire [31:0] R5690;
  wire [31:0] R5689;
  wire [31:0] R5688;
  wire [31:0] R5687;
  wire [31:0] R5686;
  wire [31:0] R5685;
  wire [31:0] R5684;
  wire [31:0] R5683;
  wire [31:0] R5682;
  wire [31:0] R5681;
  wire [31:0] R5680;
  wire [31:0] R5679;
  wire [31:0] R5678;
  wire [31:0] R5677;
  wire [31:0] R5676;
  wire [31:0] R5675;
  wire [31:0] R5674;
  wire [31:0] R5673;
  wire [31:0] R5672;
  wire [31:0] R5671;
  wire [31:0] R5670;
  wire [31:0] R5669;
  wire [31:0] R5668;
  wire [31:0] R5667;
  wire [31:0] R5666;
  wire [31:0] R5665;
  wire [31:0] R5664;
  wire [31:0] R5663;
  wire [31:0] R5662;
  wire [31:0] R5661;
  wire [31:0] R5660;
  wire [31:0] R5659;
  wire [31:0] R5658;
  wire [31:0] R5657;
  wire [31:0] R5656;
  wire [31:0] R5655;
  wire [31:0] R5654;
  wire [31:0] R5653;
  wire [31:0] R5652;
  wire [31:0] R5651;
  wire [31:0] R5650;
  wire [31:0] R5649;
  wire [31:0] R5648;
  wire [31:0] R5647;
  wire [31:0] R5646;
  wire [31:0] R5645;
  wire [31:0] R5644;
  wire [31:0] R5643;
  wire [31:0] R5642;
  wire [31:0] R5641;
  wire [31:0] R5640;
  wire [31:0] R5639;
  wire [31:0] R5638;
  wire [31:0] R5637;
  wire [31:0] R5636;
  wire [31:0] R5635;
  wire [31:0] R5634;
  wire [31:0] R5633;
  wire [31:0] R5632;
  wire [31:0] R5631;
  wire [31:0] R5630;
  wire [31:0] R5629;
  wire [31:0] R5628;
  wire [31:0] R5627;
  wire [31:0] R5626;
  wire [31:0] R5625;
  wire [31:0] R5624;
  wire [31:0] R5623;
  wire [31:0] R5622;
  wire [31:0] R5621;
  wire [31:0] R5620;
  wire [31:0] R5619;
  wire [31:0] R5618;
  wire [31:0] R5617;
  wire [31:0] R5616;
  wire [31:0] R5615;
  wire [31:0] R5614;
  wire [31:0] R5613;
  wire [31:0] R5612;
  wire [31:0] R5611;
  wire [31:0] R5610;
  wire [31:0] R5609;
  wire [31:0] R5608;
  wire [31:0] R5607;
  wire [31:0] R5606;
  wire [31:0] R5605;
  wire [31:0] R5604;
  wire [31:0] R5603;
  wire [31:0] R5602;
  wire [31:0] R5601;
  wire [31:0] R5600;
  wire [31:0] R5599;
  wire [31:0] R5598;
  wire [31:0] R5597;
  wire [31:0] R5596;
  wire [31:0] R5595;
  wire [31:0] R5594;
  wire [63:0] R5593;
  wire [31:0] R5592;
  wire [31:0] R5591;
  wire [63:0] R5590;
  wire [31:0] R5589;
  wire [63:0] R5588;
  wire [63:0] R5587;
  wire [63:0] R5586;
  wire [63:0] R5585;
  wire [63:0] R5584;
  wire [63:0] R5583;
  wire [31:0] R5582;
  wire [63:0] R5581;
  wire [63:0] R5580;
  wire [63:0] R5579;
  wire [63:0] R5578;
  wire [63:0] R5577;
  wire [63:0] R5576;
  wire [63:0] R5575;
  wire [31:0] R5574;
  wire [31:0] R5573;
  wire [31:0] R5572;
  wire [63:0] R5571;
  wire [63:0] R5570;
  wire [63:0] R5569;
  wire [63:0] R5568;
  wire [63:0] R5567;
  wire [63:0] R5566;
  wire [63:0] R5565;
  wire [63:0] R5564;
  wire [63:0] R5563;
  wire [63:0] R5562;
  wire [63:0] R5561;
  wire [63:0] R5560;
  wire [63:0] R5559;
  wire [63:0] R5558;
  wire [63:0] R5557;
  wire [63:0] R5556;
  wire [63:0] R5555;
  wire [63:0] R5554;
  wire [63:0] R5553;
  wire [63:0] R5552;
  wire [63:0] R5551;
  wire [63:0] R5550;
  wire [63:0] R5549;
  wire [63:0] R5548;
  wire [0:0] R5547;
  wire [0:0] R5546;
  wire [0:0] R5545;
  wire [0:0] R5544;
  wire [0:0] R5543;
  wire [0:0] R5542;
  wire [0:0] R5541;
  wire [0:0] R5540;
  wire [0:0] R5539;
  wire [0:0] R5538;
  wire [0:0] R5537;
  wire [0:0] R5536;
  wire [0:0] R5535;
  wire [0:0] R5534;
  wire [0:0] R5533;
  wire [0:0] R5532;
  wire [0:0] R5531;
  wire [0:0] R5530;
  wire [0:0] R5529;
  wire [0:0] R5528;
  wire [0:0] R5527;
  wire [0:0] R5526;
  wire [0:0] R5525;
  wire [0:0] R5524;
  wire [0:0] R5523;
  wire [0:0] R5522;
  wire [0:0] R5521;
  wire [0:0] R5520;
  wire [0:0] R5519;
  wire [0:0] R5518;
  wire [0:0] R5517;
  wire [0:0] R5516;
  wire [0:0] R5515;
  wire [0:0] R5514;
  wire [0:0] R5513;
  wire [0:0] R5512;
  wire [0:0] R5511;
  wire [0:0] R5510;
  wire [0:0] R5509;
  wire [0:0] R5508;
  wire [0:0] R5507;
  wire [0:0] R5506;
  wire [0:0] R5505;
  wire [0:0] R5504;
  wire [0:0] R5503;
  wire [0:0] R5502;
  wire [0:0] R5501;
  wire [0:0] R5500;
  wire [0:0] R5499;
  wire [0:0] R5498;
  wire [0:0] R5497;
  wire [0:0] R5496;
  wire [0:0] R5495;
  wire [0:0] R5494;
  wire [0:0] R5493;
  wire [0:0] R5492;
  wire [0:0] R5491;
  wire [0:0] R5490;
  wire [0:0] R5489;
  wire [0:0] R5488;
  wire [0:0] R5487;
  wire [0:0] R5486;
  wire [0:0] R5485;
  wire [0:0] R5484;
  wire [0:0] R5483;
  wire [0:0] R5482;
  wire [0:0] R5481;
  wire [0:0] R5480;
  wire [0:0] R5479;
  wire [0:0] R5478;
  wire [0:0] R5477;
  wire [0:0] R5476;
  wire [0:0] R5475;
  wire [0:0] R5474;
  wire [0:0] R5473;
  wire [0:0] R5472;
  wire [0:0] R5471;
  wire [0:0] R5470;
  wire [0:0] R5469;
  wire [0:0] R5468;
  wire [0:0] R5467;
  wire [0:0] R5466;
  wire [0:0] R5465;
  wire [0:0] R5464;
  wire [0:0] R5463;
  wire [0:0] R5462;
  wire [0:0] R5461;
  wire [0:0] R5460;
  wire [0:0] R5459;
  wire [0:0] R5458;
  wire [0:0] R5457;
  wire [0:0] R5456;
  wire [0:0] R5455;
  wire [0:0] R5454;
  wire [0:0] R5453;
  wire [0:0] R5452;
  wire [0:0] R5451;
  wire [0:0] R5450;
  wire [0:0] R5449;
  wire [0:0] R5448;
  wire [0:0] R5447;
  wire [0:0] R5446;
  wire [0:0] R5445;
  wire [0:0] R5444;
  wire [0:0] R5443;
  wire [0:0] R5442;
  wire [0:0] R5441;
  wire [0:0] R5440;
  wire [0:0] R5439;
  wire [0:0] R5438;
  wire [0:0] R5437;
  wire [0:0] R5436;
  wire [0:0] R5435;
  wire [0:0] R5434;
  wire [0:0] R5433;
  wire [0:0] R5432;
  wire [0:0] R5431;
  wire [0:0] R5430;
  wire [0:0] R5429;
  wire [0:0] R5428;
  wire [0:0] R5427;
  wire [0:0] R5426;
  wire [0:0] R5425;
  wire [0:0] R5424;
  wire [0:0] R5423;
  wire [0:0] R5422;
  wire [0:0] R5421;
  wire [0:0] R5420;
  wire [0:0] R5419;
  wire [0:0] R5418;
  wire [0:0] R5417;
  wire [0:0] R5416;
  wire [0:0] R5415;
  wire [0:0] R5414;
  wire [0:0] R5413;
  wire [0:0] R5412;
  wire [0:0] R5411;
  wire [0:0] R5410;
  wire [0:0] R5409;
  wire [0:0] R5408;
  wire [0:0] R5407;
  wire [0:0] R5406;
  wire [0:0] R5405;
  wire [0:0] R5404;
  wire [0:0] R5403;
  wire [0:0] R5402;
  wire [0:0] R5401;
  wire [0:0] R5400;
  wire [0:0] R5399;
  wire [0:0] R5398;
  wire [0:0] R5397;
  wire [0:0] R5396;
  wire [63:0] R5395;
  wire [31:0] R5394;
  wire [31:0] R5393;
  wire [31:0] R5392;
  wire [31:0] R5391;
  wire [31:0] R5390;
  wire [31:0] R5389;
  wire [31:0] R5388;
  wire [31:0] R5387;
  wire [31:0] R5386;
  wire [31:0] R5385;
  wire [31:0] R5384;
  wire [31:0] R5383;
  wire [31:0] R5382;
  wire [31:0] R5381;
  wire [31:0] R5380;
  wire [31:0] R5379;
  wire [31:0] R5378;
  wire [31:0] R5377;
  wire [31:0] R5376;
  wire [31:0] R5375;
  wire [31:0] R5374;
  wire [31:0] R5373;
  wire [31:0] R5372;
  wire [31:0] R5371;
  wire [31:0] R5370;
  wire [31:0] R5369;
  wire [31:0] R5368;
  wire [31:0] R5367;
  wire [31:0] R5366;
  wire [31:0] R5365;
  wire [31:0] R5364;
  wire [31:0] R5363;
  wire [31:0] R5362;
  wire [31:0] R5361;
  wire [31:0] R5360;
  wire [31:0] R5359;
  wire [31:0] R5358;
  wire [31:0] R5357;
  wire [31:0] R5356;
  wire [31:0] R5355;
  wire [31:0] R5354;
  wire [31:0] R5353;
  wire [31:0] R5352;
  wire [31:0] R5351;
  wire [31:0] R5350;
  wire [31:0] R5349;
  wire [31:0] R5348;
  wire [31:0] R5347;
  wire [31:0] R5346;
  wire [31:0] R5345;
  wire [31:0] R5344;
  wire [31:0] R5343;
  wire [31:0] R5342;
  wire [31:0] R5341;
  wire [31:0] R5340;
  wire [31:0] R5339;
  wire [31:0] R5338;
  wire [31:0] R5337;
  wire [31:0] R5336;
  wire [31:0] R5335;
  wire [31:0] R5334;
  wire [31:0] R5333;
  wire [31:0] R5332;
  wire [31:0] R5331;
  wire [31:0] R5330;
  wire [31:0] R5329;
  wire [31:0] R5328;
  wire [31:0] R5327;
  wire [31:0] R5326;
  wire [31:0] R5325;
  wire [31:0] R5324;
  wire [31:0] R5323;
  wire [31:0] R5322;
  wire [31:0] R5321;
  wire [31:0] R5320;
  wire [31:0] R5319;
  wire [31:0] R5318;
  wire [31:0] R5317;
  wire [31:0] R5316;
  wire [31:0] R5315;
  wire [31:0] R5314;
  wire [31:0] R5313;
  wire [31:0] R5312;
  wire [31:0] R5311;
  wire [31:0] R5310;
  wire [31:0] R5309;
  wire [31:0] R5308;
  wire [31:0] R5307;
  wire [31:0] R5306;
  wire [31:0] R5305;
  wire [31:0] R5304;
  wire [31:0] R5303;
  wire [31:0] R5302;
  wire [31:0] R5301;
  wire [31:0] R5300;
  wire [31:0] R5299;
  wire [31:0] R5298;
  wire [31:0] R5297;
  wire [31:0] R5296;
  wire [31:0] R5295;
  wire [31:0] R5294;
  wire [31:0] R5293;
  wire [31:0] R5292;
  wire [31:0] R5291;
  wire [31:0] R5290;
  wire [31:0] R5289;
  wire [31:0] R5288;
  wire [31:0] R5287;
  wire [31:0] R5286;
  wire [31:0] R5285;
  wire [31:0] R5284;
  wire [31:0] R5283;
  wire [31:0] R5282;
  wire [31:0] R5281;
  wire [31:0] R5280;
  wire [31:0] R5279;
  wire [31:0] R5278;
  wire [31:0] R5277;
  wire [31:0] R5276;
  wire [31:0] R5275;
  wire [31:0] R5274;
  wire [31:0] R5273;
  wire [31:0] R5272;
  wire [31:0] R5271;
  wire [31:0] R5270;
  wire [31:0] R5269;
  wire [31:0] R5268;
  wire [31:0] R5267;
  wire [31:0] R5266;
  wire [31:0] R5265;
  wire [31:0] R5264;
  wire [31:0] R5263;
  wire [31:0] R5262;
  wire [31:0] R5261;
  wire [31:0] R5260;
  wire [31:0] R5259;
  wire [31:0] R5258;
  wire [31:0] R5257;
  wire [31:0] R5256;
  wire [31:0] R5255;
  wire [31:0] R5254;
  wire [31:0] R5253;
  wire [31:0] R5252;
  wire [31:0] R5251;
  wire [31:0] R5250;
  wire [31:0] R5249;
  wire [63:0] R5248;
  wire [63:0] R5247;
  wire [63:0] R5246;
  wire [31:0] R5245;
  wire [31:0] R5244;
  wire [31:0] R5243;
  wire [31:0] R5242;
  wire [31:0] R5241;
  wire [31:0] R5240;
  wire [31:0] R5239;
  wire [31:0] R5238;
  wire [31:0] R5237;
  wire [31:0] R5236;
  wire [31:0] R5235;
  wire [31:0] R5234;
  wire [31:0] R5233;
  wire [31:0] R5232;
  wire [31:0] R5231;
  wire [31:0] R5230;
  wire [31:0] R5229;
  wire [31:0] R5228;
  wire [31:0] R5227;
  wire [31:0] R5226;
  wire [31:0] R5225;
  wire [31:0] R5224;
  wire [31:0] R5223;
  wire [31:0] R5222;
  wire [31:0] R5221;
  wire [31:0] R5220;
  wire [31:0] R5219;
  wire [31:0] R5218;
  wire [31:0] R5217;
  wire [31:0] R5216;
  wire [31:0] R5215;
  wire [31:0] R5214;
  wire [31:0] R5213;
  wire [31:0] R5212;
  wire [31:0] R5211;
  wire [31:0] R5210;
  wire [31:0] R5209;
  wire [31:0] R5208;
  wire [31:0] R5207;
  wire [31:0] R5206;
  wire [31:0] R5205;
  wire [31:0] R5204;
  wire [31:0] R5203;
  wire [31:0] R5202;
  wire [31:0] R5201;
  wire [31:0] R5200;
  wire [31:0] R5199;
  wire [31:0] R5198;
  wire [31:0] R5197;
  wire [31:0] R5196;
  wire [31:0] R5195;
  wire [31:0] R5194;
  wire [31:0] R5193;
  wire [31:0] R5192;
  wire [31:0] R5191;
  wire [31:0] R5190;
  wire [31:0] R5189;
  wire [31:0] R5188;
  wire [31:0] R5187;
  wire [31:0] R5186;
  wire [31:0] R5185;
  wire [31:0] R5184;
  wire [31:0] R5183;
  wire [31:0] R5182;
  wire [31:0] R5181;
  wire [31:0] R5180;
  wire [31:0] R5179;
  wire [31:0] R5178;
  wire [31:0] R5177;
  wire [31:0] R5176;
  wire [31:0] R5175;
  wire [31:0] R5174;
  wire [31:0] R5173;
  wire [31:0] R5172;
  wire [31:0] R5171;
  wire [31:0] R5170;
  wire [31:0] R5169;
  wire [31:0] R5168;
  wire [31:0] R5167;
  wire [31:0] R5166;
  wire [31:0] R5165;
  wire [31:0] R5164;
  wire [31:0] R5163;
  wire [31:0] R5162;
  wire [31:0] R5161;
  wire [31:0] R5160;
  wire [31:0] R5159;
  wire [31:0] R5158;
  wire [31:0] R5157;
  wire [31:0] R5156;
  wire [31:0] R5155;
  wire [31:0] R5154;
  wire [31:0] R5153;
  wire [31:0] R5152;
  wire [31:0] R5151;
  wire [31:0] R5150;
  wire [31:0] R5149;
  wire [31:0] R5148;
  wire [31:0] R5147;
  wire [31:0] R5146;
  wire [31:0] R5145;
  wire [31:0] R5144;
  wire [31:0] R5143;
  wire [31:0] R5142;
  wire [31:0] R5141;
  wire [31:0] R5140;
  wire [31:0] R5139;
  wire [31:0] R5138;
  wire [31:0] R5137;
  wire [31:0] R5136;
  wire [31:0] R5135;
  wire [31:0] R5134;
  wire [31:0] R5133;
  wire [31:0] R5132;
  wire [31:0] R5131;
  wire [31:0] R5130;
  wire [31:0] R5129;
  wire [31:0] R5128;
  wire [31:0] R5127;
  wire [31:0] R5126;
  wire [31:0] R5125;
  wire [31:0] R5124;
  wire [31:0] R5123;
  wire [31:0] R5122;
  wire [31:0] R5121;
  wire [31:0] R5120;
  wire [31:0] R5119;
  wire [31:0] R5118;
  wire [31:0] R5117;
  wire [31:0] R5116;
  wire [31:0] R5115;
  wire [31:0] R5114;
  wire [31:0] R5113;
  wire [31:0] R5112;
  wire [31:0] R5111;
  wire [31:0] R5110;
  wire [31:0] R5109;
  wire [31:0] R5108;
  wire [31:0] R5107;
  wire [31:0] R5106;
  wire [31:0] R5105;
  wire [31:0] R5104;
  wire [31:0] R5103;
  wire [31:0] R5102;
  wire [31:0] R5101;
  wire [31:0] R5100;
  wire [31:0] R5099;
  wire [31:0] R5098;
  wire [31:0] R5097;
  wire [31:0] R5096;
  wire [31:0] R5095;
  wire [31:0] R5094;
  wire [31:0] R5093;
  wire [63:0] R5092;
  wire [31:0] R5091;
  wire [31:0] R5090;
  wire [63:0] R5089;
  wire [31:0] R5088;
  wire [63:0] R5087;
  wire [63:0] R5086;
  wire [63:0] R5085;
  wire [63:0] R5084;
  wire [63:0] R5083;
  wire [63:0] R5082;
  wire [31:0] R5081;
  wire [63:0] R5080;
  wire [63:0] R5079;
  wire [63:0] R5078;
  wire [63:0] R5077;
  wire [63:0] R5076;
  wire [63:0] R5075;
  wire [63:0] R5074;
  wire [31:0] R5073;
  wire [31:0] R5072;
  wire [31:0] R5071;
  wire [63:0] R5070;
  wire [63:0] R5069;
  wire [63:0] R5068;
  wire [63:0] R5067;
  wire [63:0] R5066;
  wire [63:0] R5065;
  wire [63:0] R5064;
  wire [63:0] R5063;
  wire [63:0] R5062;
  wire [63:0] R5061;
  wire [63:0] R5060;
  wire [63:0] R5059;
  wire [63:0] R5058;
  wire [63:0] R5057;
  wire [63:0] R5056;
  wire [63:0] R5055;
  wire [63:0] R5054;
  wire [63:0] R5053;
  wire [63:0] R5052;
  wire [63:0] R5051;
  wire [63:0] R5050;
  wire [63:0] R5049;
  wire [63:0] R5048;
  wire [63:0] R5047;
  wire [0:0] R5046;
  wire [0:0] R5045;
  wire [0:0] R5044;
  wire [0:0] R5043;
  wire [0:0] R5042;
  wire [0:0] R5041;
  wire [0:0] R5040;
  wire [0:0] R5039;
  wire [0:0] R5038;
  wire [0:0] R5037;
  wire [0:0] R5036;
  wire [0:0] R5035;
  wire [0:0] R5034;
  wire [0:0] R5033;
  wire [0:0] R5032;
  wire [0:0] R5031;
  wire [0:0] R5030;
  wire [0:0] R5029;
  wire [0:0] R5028;
  wire [0:0] R5027;
  wire [0:0] R5026;
  wire [0:0] R5025;
  wire [0:0] R5024;
  wire [0:0] R5023;
  wire [0:0] R5022;
  wire [0:0] R5021;
  wire [0:0] R5020;
  wire [0:0] R5019;
  wire [0:0] R5018;
  wire [0:0] R5017;
  wire [0:0] R5016;
  wire [0:0] R5015;
  wire [0:0] R5014;
  wire [0:0] R5013;
  wire [0:0] R5012;
  wire [0:0] R5011;
  wire [0:0] R5010;
  wire [0:0] R5009;
  wire [0:0] R5008;
  wire [0:0] R5007;
  wire [0:0] R5006;
  wire [0:0] R5005;
  wire [0:0] R5004;
  wire [0:0] R5003;
  wire [0:0] R5002;
  wire [0:0] R5001;
  wire [0:0] R5000;
  wire [0:0] R4999;
  wire [0:0] R4998;
  wire [0:0] R4997;
  wire [0:0] R4996;
  wire [0:0] R4995;
  wire [0:0] R4994;
  wire [0:0] R4993;
  wire [0:0] R4992;
  wire [0:0] R4991;
  wire [0:0] R4990;
  wire [0:0] R4989;
  wire [0:0] R4988;
  wire [0:0] R4987;
  wire [0:0] R4986;
  wire [0:0] R4985;
  wire [0:0] R4984;
  wire [0:0] R4983;
  wire [0:0] R4982;
  wire [0:0] R4981;
  wire [0:0] R4980;
  wire [0:0] R4979;
  wire [0:0] R4978;
  wire [0:0] R4977;
  wire [0:0] R4976;
  wire [0:0] R4975;
  wire [0:0] R4974;
  wire [0:0] R4973;
  wire [0:0] R4972;
  wire [0:0] R4971;
  wire [0:0] R4970;
  wire [0:0] R4969;
  wire [0:0] R4968;
  wire [0:0] R4967;
  wire [0:0] R4966;
  wire [0:0] R4965;
  wire [0:0] R4964;
  wire [0:0] R4963;
  wire [0:0] R4962;
  wire [0:0] R4961;
  wire [0:0] R4960;
  wire [0:0] R4959;
  wire [0:0] R4958;
  wire [0:0] R4957;
  wire [0:0] R4956;
  wire [0:0] R4955;
  wire [0:0] R4954;
  wire [0:0] R4953;
  wire [0:0] R4952;
  wire [0:0] R4951;
  wire [0:0] R4950;
  wire [0:0] R4949;
  wire [0:0] R4948;
  wire [0:0] R4947;
  wire [0:0] R4946;
  wire [0:0] R4945;
  wire [0:0] R4944;
  wire [0:0] R4943;
  wire [0:0] R4942;
  wire [0:0] R4941;
  wire [0:0] R4940;
  wire [0:0] R4939;
  wire [0:0] R4938;
  wire [0:0] R4937;
  wire [0:0] R4936;
  wire [0:0] R4935;
  wire [0:0] R4934;
  wire [0:0] R4933;
  wire [0:0] R4932;
  wire [0:0] R4931;
  wire [0:0] R4930;
  wire [0:0] R4929;
  wire [0:0] R4928;
  wire [0:0] R4927;
  wire [0:0] R4926;
  wire [0:0] R4925;
  wire [0:0] R4924;
  wire [0:0] R4923;
  wire [0:0] R4922;
  wire [0:0] R4921;
  wire [0:0] R4920;
  wire [0:0] R4919;
  wire [0:0] R4918;
  wire [0:0] R4917;
  wire [0:0] R4916;
  wire [0:0] R4915;
  wire [0:0] R4914;
  wire [0:0] R4913;
  wire [0:0] R4912;
  wire [0:0] R4911;
  wire [0:0] R4910;
  wire [0:0] R4909;
  wire [0:0] R4908;
  wire [0:0] R4907;
  wire [0:0] R4906;
  wire [0:0] R4905;
  wire [0:0] R4904;
  wire [0:0] R4903;
  wire [0:0] R4902;
  wire [0:0] R4901;
  wire [0:0] R4900;
  wire [0:0] R4899;
  wire [0:0] R4898;
  wire [0:0] R4897;
  wire [0:0] R4896;
  wire [0:0] R4895;
  wire [0:0] R4894;
  wire [0:0] R4893;
  wire [0:0] R4892;
  wire [0:0] R4891;
  wire [0:0] R4890;
  wire [0:0] R4889;
  wire [0:0] R4888;
  wire [0:0] R4887;
  wire [0:0] R4886;
  wire [0:0] R4885;
  wire [0:0] R4884;
  wire [0:0] R4883;
  wire [0:0] R4882;
  wire [0:0] R4881;
  wire [63:0] R4880;
  wire [31:0] R4879;
  wire [31:0] R4878;
  wire [31:0] R4877;
  wire [31:0] R4876;
  wire [31:0] R4875;
  wire [31:0] R4874;
  wire [31:0] R4873;
  wire [31:0] R4872;
  wire [31:0] R4871;
  wire [31:0] R4870;
  wire [31:0] R4869;
  wire [31:0] R4868;
  wire [31:0] R4867;
  wire [31:0] R4866;
  wire [31:0] R4865;
  wire [31:0] R4864;
  wire [31:0] R4863;
  wire [31:0] R4862;
  wire [31:0] R4861;
  wire [31:0] R4860;
  wire [31:0] R4859;
  wire [31:0] R4858;
  wire [31:0] R4857;
  wire [31:0] R4856;
  wire [31:0] R4855;
  wire [31:0] R4854;
  wire [31:0] R4853;
  wire [31:0] R4852;
  wire [31:0] R4851;
  wire [31:0] R4850;
  wire [31:0] R4849;
  wire [31:0] R4848;
  wire [31:0] R4847;
  wire [31:0] R4846;
  wire [31:0] R4845;
  wire [31:0] R4844;
  wire [31:0] R4843;
  wire [31:0] R4842;
  wire [31:0] R4841;
  wire [31:0] R4840;
  wire [31:0] R4839;
  wire [31:0] R4838;
  wire [31:0] R4837;
  wire [31:0] R4836;
  wire [31:0] R4835;
  wire [31:0] R4834;
  wire [31:0] R4833;
  wire [31:0] R4832;
  wire [31:0] R4831;
  wire [31:0] R4830;
  wire [31:0] R4829;
  wire [31:0] R4828;
  wire [31:0] R4827;
  wire [31:0] R4826;
  wire [31:0] R4825;
  wire [31:0] R4824;
  wire [31:0] R4823;
  wire [31:0] R4822;
  wire [31:0] R4821;
  wire [31:0] R4820;
  wire [31:0] R4819;
  wire [31:0] R4818;
  wire [31:0] R4817;
  wire [31:0] R4816;
  wire [31:0] R4815;
  wire [31:0] R4814;
  wire [31:0] R4813;
  wire [31:0] R4812;
  wire [31:0] R4811;
  wire [31:0] R4810;
  wire [31:0] R4809;
  wire [31:0] R4808;
  wire [31:0] R4807;
  wire [31:0] R4806;
  wire [31:0] R4805;
  wire [31:0] R4804;
  wire [31:0] R4803;
  wire [31:0] R4802;
  wire [31:0] R4801;
  wire [31:0] R4800;
  wire [31:0] R4799;
  wire [31:0] R4798;
  wire [31:0] R4797;
  wire [31:0] R4796;
  wire [31:0] R4795;
  wire [31:0] R4794;
  wire [31:0] R4793;
  wire [31:0] R4792;
  wire [31:0] R4791;
  wire [31:0] R4790;
  wire [31:0] R4789;
  wire [31:0] R4788;
  wire [31:0] R4787;
  wire [31:0] R4786;
  wire [31:0] R4785;
  wire [31:0] R4784;
  wire [31:0] R4783;
  wire [31:0] R4782;
  wire [31:0] R4781;
  wire [31:0] R4780;
  wire [31:0] R4779;
  wire [31:0] R4778;
  wire [31:0] R4777;
  wire [31:0] R4776;
  wire [31:0] R4775;
  wire [31:0] R4774;
  wire [31:0] R4773;
  wire [31:0] R4772;
  wire [31:0] R4771;
  wire [31:0] R4770;
  wire [31:0] R4769;
  wire [31:0] R4768;
  wire [31:0] R4767;
  wire [31:0] R4766;
  wire [31:0] R4765;
  wire [31:0] R4764;
  wire [31:0] R4763;
  wire [31:0] R4762;
  wire [31:0] R4761;
  wire [31:0] R4760;
  wire [31:0] R4759;
  wire [31:0] R4758;
  wire [31:0] R4757;
  wire [31:0] R4756;
  wire [31:0] R4755;
  wire [31:0] R4754;
  wire [31:0] R4753;
  wire [31:0] R4752;
  wire [31:0] R4751;
  wire [31:0] R4750;
  wire [31:0] R4749;
  wire [31:0] R4748;
  wire [31:0] R4747;
  wire [31:0] R4746;
  wire [31:0] R4745;
  wire [31:0] R4744;
  wire [31:0] R4743;
  wire [31:0] R4742;
  wire [31:0] R4741;
  wire [31:0] R4740;
  wire [31:0] R4739;
  wire [31:0] R4738;
  wire [31:0] R4737;
  wire [31:0] R4736;
  wire [31:0] R4735;
  wire [31:0] R4734;
  wire [31:0] R4733;
  wire [31:0] R4732;
  wire [31:0] R4731;
  wire [31:0] R4730;
  wire [31:0] R4729;
  wire [31:0] R4728;
  wire [31:0] R4727;
  wire [31:0] R4726;
  wire [31:0] R4725;
  wire [31:0] R4724;
  wire [31:0] R4723;
  wire [31:0] R4722;
  wire [31:0] R4721;
  wire [31:0] R4720;
  wire [63:0] R4719;
  wire [63:0] R4718;
  wire [63:0] R4717;
  wire [31:0] R4716;
  wire [31:0] R4715;
  wire [31:0] R4714;
  wire [31:0] R4713;
  wire [31:0] R4712;
  wire [31:0] R4711;
  wire [31:0] R4710;
  wire [31:0] R4709;
  wire [31:0] R4708;
  wire [31:0] R4707;
  wire [31:0] R4706;
  wire [31:0] R4705;
  wire [31:0] R4704;
  wire [31:0] R4703;
  wire [31:0] R4702;
  wire [31:0] R4701;
  wire [31:0] R4700;
  wire [31:0] R4699;
  wire [31:0] R4698;
  wire [31:0] R4697;
  wire [31:0] R4696;
  wire [31:0] R4695;
  wire [31:0] R4694;
  wire [31:0] R4693;
  wire [31:0] R4692;
  wire [31:0] R4691;
  wire [31:0] R4690;
  wire [31:0] R4689;
  wire [31:0] R4688;
  wire [31:0] R4687;
  wire [31:0] R4686;
  wire [31:0] R4685;
  wire [31:0] R4684;
  wire [31:0] R4683;
  wire [31:0] R4682;
  wire [31:0] R4681;
  wire [31:0] R4680;
  wire [31:0] R4679;
  wire [31:0] R4678;
  wire [31:0] R4677;
  wire [31:0] R4676;
  wire [31:0] R4675;
  wire [31:0] R4674;
  wire [31:0] R4673;
  wire [31:0] R4672;
  wire [31:0] R4671;
  wire [31:0] R4670;
  wire [31:0] R4669;
  wire [31:0] R4668;
  wire [31:0] R4667;
  wire [31:0] R4666;
  wire [31:0] R4665;
  wire [31:0] R4664;
  wire [31:0] R4663;
  wire [31:0] R4662;
  wire [31:0] R4661;
  wire [31:0] R4660;
  wire [31:0] R4659;
  wire [31:0] R4658;
  wire [31:0] R4657;
  wire [31:0] R4656;
  wire [31:0] R4655;
  wire [31:0] R4654;
  wire [31:0] R4653;
  wire [31:0] R4652;
  wire [31:0] R4651;
  wire [31:0] R4650;
  wire [31:0] R4649;
  wire [31:0] R4648;
  wire [31:0] R4647;
  wire [31:0] R4646;
  wire [31:0] R4645;
  wire [31:0] R4644;
  wire [31:0] R4643;
  wire [31:0] R4642;
  wire [31:0] R4641;
  wire [31:0] R4640;
  wire [31:0] R4639;
  wire [31:0] R4638;
  wire [31:0] R4637;
  wire [31:0] R4636;
  wire [31:0] R4635;
  wire [31:0] R4634;
  wire [31:0] R4633;
  wire [31:0] R4632;
  wire [31:0] R4631;
  wire [31:0] R4630;
  wire [31:0] R4629;
  wire [31:0] R4628;
  wire [31:0] R4627;
  wire [31:0] R4626;
  wire [31:0] R4625;
  wire [31:0] R4624;
  wire [31:0] R4623;
  wire [31:0] R4622;
  wire [31:0] R4621;
  wire [31:0] R4620;
  wire [31:0] R4619;
  wire [31:0] R4618;
  wire [31:0] R4617;
  wire [31:0] R4616;
  wire [31:0] R4615;
  wire [31:0] R4614;
  wire [31:0] R4613;
  wire [31:0] R4612;
  wire [31:0] R4611;
  wire [31:0] R4610;
  wire [31:0] R4609;
  wire [31:0] R4608;
  wire [31:0] R4607;
  wire [31:0] R4606;
  wire [31:0] R4605;
  wire [31:0] R4604;
  wire [31:0] R4603;
  wire [31:0] R4602;
  wire [31:0] R4601;
  wire [31:0] R4600;
  wire [31:0] R4599;
  wire [31:0] R4598;
  wire [31:0] R4597;
  wire [31:0] R4596;
  wire [31:0] R4595;
  wire [31:0] R4594;
  wire [31:0] R4593;
  wire [31:0] R4592;
  wire [31:0] R4591;
  wire [31:0] R4590;
  wire [31:0] R4589;
  wire [31:0] R4588;
  wire [31:0] R4587;
  wire [31:0] R4586;
  wire [31:0] R4585;
  wire [31:0] R4584;
  wire [31:0] R4583;
  wire [31:0] R4582;
  wire [31:0] R4581;
  wire [31:0] R4580;
  wire [31:0] R4579;
  wire [31:0] R4578;
  wire [31:0] R4577;
  wire [31:0] R4576;
  wire [31:0] R4575;
  wire [31:0] R4574;
  wire [31:0] R4573;
  wire [31:0] R4572;
  wire [31:0] R4571;
  wire [31:0] R4570;
  wire [31:0] R4569;
  wire [31:0] R4568;
  wire [31:0] R4567;
  wire [31:0] R4566;
  wire [31:0] R4565;
  wire [31:0] R4564;
  wire [31:0] R4563;
  wire [31:0] R4562;
  wire [31:0] R4561;
  wire [31:0] R4560;
  wire [31:0] R4559;
  wire [31:0] R4558;
  wire [31:0] R4557;
  wire [31:0] R4556;
  wire [31:0] R4555;
  wire [31:0] R4554;
  wire [31:0] R4553;
  wire [31:0] R4552;
  wire [31:0] R4551;
  wire [31:0] R4550;
  wire [63:0] R4549;
  wire [31:0] R4548;
  wire [31:0] R4547;
  wire [63:0] R4546;
  wire [31:0] R4545;
  wire [63:0] R4544;
  wire [63:0] R4543;
  wire [63:0] R4542;
  wire [63:0] R4541;
  wire [63:0] R4540;
  wire [63:0] R4539;
  wire [31:0] R4538;
  wire [63:0] R4537;
  wire [63:0] R4536;
  wire [63:0] R4535;
  wire [63:0] R4534;
  wire [63:0] R4533;
  wire [63:0] R4532;
  wire [63:0] R4531;
  wire [31:0] R4530;
  wire [31:0] R4529;
  wire [31:0] R4528;
  wire [63:0] R4527;
  wire [63:0] R4526;
  wire [63:0] R4525;
  wire [63:0] R4524;
  wire [63:0] R4523;
  wire [63:0] R4522;
  wire [63:0] R4521;
  wire [63:0] R4520;
  wire [63:0] R4519;
  wire [63:0] R4518;
  wire [63:0] R4517;
  wire [63:0] R4516;
  wire [63:0] R4515;
  wire [63:0] R4514;
  wire [63:0] R4513;
  wire [63:0] R4512;
  wire [63:0] R4511;
  wire [63:0] R4510;
  wire [63:0] R4509;
  wire [63:0] R4508;
  wire [63:0] R4507;
  wire [63:0] R4506;
  wire [63:0] R4505;
  wire [63:0] R4504;
  wire [0:0] R4503;
  wire [0:0] R4502;
  wire [0:0] R4501;
  wire [0:0] R4500;
  wire [0:0] R4499;
  wire [0:0] R4498;
  wire [0:0] R4497;
  wire [0:0] R4496;
  wire [0:0] R4495;
  wire [0:0] R4494;
  wire [0:0] R4493;
  wire [0:0] R4492;
  wire [0:0] R4491;
  wire [0:0] R4490;
  wire [0:0] R4489;
  wire [0:0] R4488;
  wire [0:0] R4487;
  wire [0:0] R4486;
  wire [0:0] R4485;
  wire [0:0] R4484;
  wire [0:0] R4483;
  wire [0:0] R4482;
  wire [0:0] R4481;
  wire [0:0] R4480;
  wire [0:0] R4479;
  wire [0:0] R4478;
  wire [0:0] R4477;
  wire [0:0] R4476;
  wire [0:0] R4475;
  wire [0:0] R4474;
  wire [0:0] R4473;
  wire [0:0] R4472;
  wire [0:0] R4471;
  wire [0:0] R4470;
  wire [0:0] R4469;
  wire [0:0] R4468;
  wire [0:0] R4467;
  wire [0:0] R4466;
  wire [0:0] R4465;
  wire [0:0] R4464;
  wire [0:0] R4463;
  wire [0:0] R4462;
  wire [0:0] R4461;
  wire [0:0] R4460;
  wire [0:0] R4459;
  wire [0:0] R4458;
  wire [0:0] R4457;
  wire [0:0] R4456;
  wire [0:0] R4455;
  wire [0:0] R4454;
  wire [0:0] R4453;
  wire [0:0] R4452;
  wire [0:0] R4451;
  wire [0:0] R4450;
  wire [0:0] R4449;
  wire [0:0] R4448;
  wire [0:0] R4447;
  wire [0:0] R4446;
  wire [0:0] R4445;
  wire [0:0] R4444;
  wire [0:0] R4443;
  wire [0:0] R4442;
  wire [0:0] R4441;
  wire [0:0] R4440;
  wire [0:0] R4439;
  wire [0:0] R4438;
  wire [0:0] R4437;
  wire [0:0] R4436;
  wire [0:0] R4435;
  wire [0:0] R4434;
  wire [0:0] R4433;
  wire [0:0] R4432;
  wire [0:0] R4431;
  wire [0:0] R4430;
  wire [0:0] R4429;
  wire [0:0] R4428;
  wire [0:0] R4427;
  wire [0:0] R4426;
  wire [0:0] R4425;
  wire [0:0] R4424;
  wire [0:0] R4423;
  wire [0:0] R4422;
  wire [0:0] R4421;
  wire [0:0] R4420;
  wire [0:0] R4419;
  wire [0:0] R4418;
  wire [0:0] R4417;
  wire [0:0] R4416;
  wire [0:0] R4415;
  wire [0:0] R4414;
  wire [0:0] R4413;
  wire [0:0] R4412;
  wire [0:0] R4411;
  wire [0:0] R4410;
  wire [0:0] R4409;
  wire [0:0] R4408;
  wire [0:0] R4407;
  wire [0:0] R4406;
  wire [0:0] R4405;
  wire [0:0] R4404;
  wire [0:0] R4403;
  wire [0:0] R4402;
  wire [0:0] R4401;
  wire [0:0] R4400;
  wire [0:0] R4399;
  wire [0:0] R4398;
  wire [0:0] R4397;
  wire [0:0] R4396;
  wire [0:0] R4395;
  wire [0:0] R4394;
  wire [0:0] R4393;
  wire [0:0] R4392;
  wire [0:0] R4391;
  wire [0:0] R4390;
  wire [0:0] R4389;
  wire [0:0] R4388;
  wire [0:0] R4387;
  wire [0:0] R4386;
  wire [0:0] R4385;
  wire [0:0] R4384;
  wire [0:0] R4383;
  wire [0:0] R4382;
  wire [0:0] R4381;
  wire [0:0] R4380;
  wire [0:0] R4379;
  wire [0:0] R4378;
  wire [0:0] R4377;
  wire [0:0] R4376;
  wire [0:0] R4375;
  wire [0:0] R4374;
  wire [0:0] R4373;
  wire [0:0] R4372;
  wire [0:0] R4371;
  wire [0:0] R4370;
  wire [0:0] R4369;
  wire [0:0] R4368;
  wire [0:0] R4367;
  wire [0:0] R4366;
  wire [0:0] R4365;
  wire [0:0] R4364;
  wire [0:0] R4363;
  wire [0:0] R4362;
  wire [0:0] R4361;
  wire [0:0] R4360;
  wire [0:0] R4359;
  wire [0:0] R4358;
  wire [0:0] R4357;
  wire [0:0] R4356;
  wire [0:0] R4355;
  wire [0:0] R4354;
  wire [0:0] R4353;
  wire [0:0] R4352;
  wire [0:0] R4351;
  wire [0:0] R4350;
  wire [0:0] R4349;
  wire [0:0] R4348;
  wire [0:0] R4347;
  wire [0:0] R4346;
  wire [0:0] R4345;
  wire [0:0] R4344;
  wire [0:0] R4343;
  wire [0:0] R4342;
  wire [0:0] R4341;
  wire [0:0] R4340;
  wire [0:0] R4339;
  wire [0:0] R4338;
  wire [0:0] R4337;
  wire [0:0] R4336;
  wire [0:0] R4335;
  wire [0:0] R4334;
  wire [0:0] R4333;
  wire [0:0] R4332;
  wire [0:0] R4331;
  wire [0:0] R4330;
  wire [0:0] R4329;
  wire [0:0] R4328;
  wire [0:0] R4327;
  wire [0:0] R4326;
  wire [0:0] R4325;
  wire [0:0] R4324;
  wire [63:0] R4323;
  wire [31:0] R4322;
  wire [31:0] R4321;
  wire [31:0] R4320;
  wire [31:0] R4319;
  wire [31:0] R4318;
  wire [31:0] R4317;
  wire [31:0] R4316;
  wire [31:0] R4315;
  wire [31:0] R4314;
  wire [31:0] R4313;
  wire [31:0] R4312;
  wire [31:0] R4311;
  wire [31:0] R4310;
  wire [31:0] R4309;
  wire [31:0] R4308;
  wire [31:0] R4307;
  wire [31:0] R4306;
  wire [31:0] R4305;
  wire [31:0] R4304;
  wire [31:0] R4303;
  wire [31:0] R4302;
  wire [31:0] R4301;
  wire [31:0] R4300;
  wire [31:0] R4299;
  wire [31:0] R4298;
  wire [31:0] R4297;
  wire [31:0] R4296;
  wire [31:0] R4295;
  wire [31:0] R4294;
  wire [31:0] R4293;
  wire [31:0] R4292;
  wire [31:0] R4291;
  wire [31:0] R4290;
  wire [31:0] R4289;
  wire [31:0] R4288;
  wire [31:0] R4287;
  wire [31:0] R4286;
  wire [31:0] R4285;
  wire [31:0] R4284;
  wire [31:0] R4283;
  wire [31:0] R4282;
  wire [31:0] R4281;
  wire [31:0] R4280;
  wire [31:0] R4279;
  wire [31:0] R4278;
  wire [31:0] R4277;
  wire [31:0] R4276;
  wire [31:0] R4275;
  wire [31:0] R4274;
  wire [31:0] R4273;
  wire [31:0] R4272;
  wire [31:0] R4271;
  wire [31:0] R4270;
  wire [31:0] R4269;
  wire [31:0] R4268;
  wire [31:0] R4267;
  wire [31:0] R4266;
  wire [31:0] R4265;
  wire [31:0] R4264;
  wire [31:0] R4263;
  wire [31:0] R4262;
  wire [31:0] R4261;
  wire [31:0] R4260;
  wire [31:0] R4259;
  wire [31:0] R4258;
  wire [31:0] R4257;
  wire [31:0] R4256;
  wire [31:0] R4255;
  wire [31:0] R4254;
  wire [31:0] R4253;
  wire [31:0] R4252;
  wire [31:0] R4251;
  wire [31:0] R4250;
  wire [31:0] R4249;
  wire [31:0] R4248;
  wire [31:0] R4247;
  wire [31:0] R4246;
  wire [31:0] R4245;
  wire [31:0] R4244;
  wire [31:0] R4243;
  wire [31:0] R4242;
  wire [31:0] R4241;
  wire [31:0] R4240;
  wire [31:0] R4239;
  wire [31:0] R4238;
  wire [31:0] R4237;
  wire [31:0] R4236;
  wire [31:0] R4235;
  wire [31:0] R4234;
  wire [31:0] R4233;
  wire [31:0] R4232;
  wire [31:0] R4231;
  wire [31:0] R4230;
  wire [31:0] R4229;
  wire [31:0] R4228;
  wire [31:0] R4227;
  wire [31:0] R4226;
  wire [31:0] R4225;
  wire [31:0] R4224;
  wire [31:0] R4223;
  wire [31:0] R4222;
  wire [31:0] R4221;
  wire [31:0] R4220;
  wire [31:0] R4219;
  wire [31:0] R4218;
  wire [31:0] R4217;
  wire [31:0] R4216;
  wire [31:0] R4215;
  wire [31:0] R4214;
  wire [31:0] R4213;
  wire [31:0] R4212;
  wire [31:0] R4211;
  wire [31:0] R4210;
  wire [31:0] R4209;
  wire [31:0] R4208;
  wire [31:0] R4207;
  wire [31:0] R4206;
  wire [31:0] R4205;
  wire [31:0] R4204;
  wire [31:0] R4203;
  wire [31:0] R4202;
  wire [31:0] R4201;
  wire [31:0] R4200;
  wire [31:0] R4199;
  wire [31:0] R4198;
  wire [31:0] R4197;
  wire [31:0] R4196;
  wire [31:0] R4195;
  wire [31:0] R4194;
  wire [31:0] R4193;
  wire [31:0] R4192;
  wire [31:0] R4191;
  wire [31:0] R4190;
  wire [31:0] R4189;
  wire [31:0] R4188;
  wire [31:0] R4187;
  wire [31:0] R4186;
  wire [31:0] R4185;
  wire [31:0] R4184;
  wire [31:0] R4183;
  wire [31:0] R4182;
  wire [31:0] R4181;
  wire [31:0] R4180;
  wire [31:0] R4179;
  wire [31:0] R4178;
  wire [31:0] R4177;
  wire [31:0] R4176;
  wire [31:0] R4175;
  wire [31:0] R4174;
  wire [31:0] R4173;
  wire [31:0] R4172;
  wire [31:0] R4171;
  wire [31:0] R4170;
  wire [31:0] R4169;
  wire [31:0] R4168;
  wire [31:0] R4167;
  wire [31:0] R4166;
  wire [31:0] R4165;
  wire [31:0] R4164;
  wire [31:0] R4163;
  wire [31:0] R4162;
  wire [31:0] R4161;
  wire [31:0] R4160;
  wire [31:0] R4159;
  wire [31:0] R4158;
  wire [31:0] R4157;
  wire [31:0] R4156;
  wire [31:0] R4155;
  wire [31:0] R4154;
  wire [31:0] R4153;
  wire [31:0] R4152;
  wire [31:0] R4151;
  wire [31:0] R4150;
  wire [31:0] R4149;
  wire [63:0] R4148;
  wire [63:0] R4147;
  wire [63:0] R4146;
  wire [31:0] R4145;
  wire [31:0] R4144;
  wire [31:0] R4143;
  wire [31:0] R4142;
  wire [31:0] R4141;
  wire [31:0] R4140;
  wire [31:0] R4139;
  wire [31:0] R4138;
  wire [31:0] R4137;
  wire [31:0] R4136;
  wire [31:0] R4135;
  wire [31:0] R4134;
  wire [31:0] R4133;
  wire [31:0] R4132;
  wire [31:0] R4131;
  wire [31:0] R4130;
  wire [31:0] R4129;
  wire [31:0] R4128;
  wire [31:0] R4127;
  wire [31:0] R4126;
  wire [31:0] R4125;
  wire [31:0] R4124;
  wire [31:0] R4123;
  wire [31:0] R4122;
  wire [31:0] R4121;
  wire [31:0] R4120;
  wire [31:0] R4119;
  wire [31:0] R4118;
  wire [31:0] R4117;
  wire [31:0] R4116;
  wire [31:0] R4115;
  wire [31:0] R4114;
  wire [31:0] R4113;
  wire [31:0] R4112;
  wire [31:0] R4111;
  wire [31:0] R4110;
  wire [31:0] R4109;
  wire [31:0] R4108;
  wire [31:0] R4107;
  wire [31:0] R4106;
  wire [31:0] R4105;
  wire [31:0] R4104;
  wire [31:0] R4103;
  wire [31:0] R4102;
  wire [31:0] R4101;
  wire [31:0] R4100;
  wire [31:0] R4099;
  wire [31:0] R4098;
  wire [31:0] R4097;
  wire [31:0] R4096;
  wire [31:0] R4095;
  wire [31:0] R4094;
  wire [31:0] R4093;
  wire [31:0] R4092;
  wire [31:0] R4091;
  wire [31:0] R4090;
  wire [31:0] R4089;
  wire [31:0] R4088;
  wire [31:0] R4087;
  wire [31:0] R4086;
  wire [31:0] R4085;
  wire [31:0] R4084;
  wire [31:0] R4083;
  wire [31:0] R4082;
  wire [31:0] R4081;
  wire [31:0] R4080;
  wire [31:0] R4079;
  wire [31:0] R4078;
  wire [31:0] R4077;
  wire [31:0] R4076;
  wire [31:0] R4075;
  wire [31:0] R4074;
  wire [31:0] R4073;
  wire [31:0] R4072;
  wire [31:0] R4071;
  wire [31:0] R4070;
  wire [31:0] R4069;
  wire [31:0] R4068;
  wire [31:0] R4067;
  wire [31:0] R4066;
  wire [31:0] R4065;
  wire [31:0] R4064;
  wire [31:0] R4063;
  wire [31:0] R4062;
  wire [31:0] R4061;
  wire [31:0] R4060;
  wire [31:0] R4059;
  wire [31:0] R4058;
  wire [31:0] R4057;
  wire [31:0] R4056;
  wire [31:0] R4055;
  wire [31:0] R4054;
  wire [31:0] R4053;
  wire [31:0] R4052;
  wire [31:0] R4051;
  wire [31:0] R4050;
  wire [31:0] R4049;
  wire [31:0] R4048;
  wire [31:0] R4047;
  wire [31:0] R4046;
  wire [31:0] R4045;
  wire [31:0] R4044;
  wire [31:0] R4043;
  wire [31:0] R4042;
  wire [31:0] R4041;
  wire [31:0] R4040;
  wire [31:0] R4039;
  wire [31:0] R4038;
  wire [31:0] R4037;
  wire [31:0] R4036;
  wire [31:0] R4035;
  wire [31:0] R4034;
  wire [31:0] R4033;
  wire [31:0] R4032;
  wire [31:0] R4031;
  wire [31:0] R4030;
  wire [31:0] R4029;
  wire [31:0] R4028;
  wire [31:0] R4027;
  wire [31:0] R4026;
  wire [31:0] R4025;
  wire [31:0] R4024;
  wire [31:0] R4023;
  wire [31:0] R4022;
  wire [31:0] R4021;
  wire [31:0] R4020;
  wire [31:0] R4019;
  wire [31:0] R4018;
  wire [31:0] R4017;
  wire [31:0] R4016;
  wire [31:0] R4015;
  wire [31:0] R4014;
  wire [31:0] R4013;
  wire [31:0] R4012;
  wire [31:0] R4011;
  wire [31:0] R4010;
  wire [31:0] R4009;
  wire [31:0] R4008;
  wire [31:0] R4007;
  wire [31:0] R4006;
  wire [31:0] R4005;
  wire [31:0] R4004;
  wire [31:0] R4003;
  wire [31:0] R4002;
  wire [31:0] R4001;
  wire [31:0] R4000;
  wire [31:0] R3999;
  wire [31:0] R3998;
  wire [31:0] R3997;
  wire [31:0] R3996;
  wire [31:0] R3995;
  wire [31:0] R3994;
  wire [31:0] R3993;
  wire [31:0] R3992;
  wire [31:0] R3991;
  wire [31:0] R3990;
  wire [31:0] R3989;
  wire [31:0] R3988;
  wire [31:0] R3987;
  wire [31:0] R3986;
  wire [31:0] R3985;
  wire [31:0] R3984;
  wire [31:0] R3983;
  wire [31:0] R3982;
  wire [31:0] R3981;
  wire [31:0] R3980;
  wire [31:0] R3979;
  wire [31:0] R3978;
  wire [31:0] R3977;
  wire [31:0] R3976;
  wire [31:0] R3975;
  wire [31:0] R3974;
  wire [31:0] R3973;
  wire [31:0] R3972;
  wire [31:0] R3971;
  wire [31:0] R3970;
  wire [31:0] R3969;
  wire [31:0] R3968;
  wire [31:0] R3967;
  wire [31:0] R3966;
  wire [31:0] R3965;
  wire [63:0] R3964;
  wire [31:0] R3963;
  wire [31:0] R3962;
  wire [63:0] R3961;
  wire [31:0] R3960;
  wire [63:0] R3959;
  wire [63:0] R3958;
  wire [63:0] R3957;
  wire [63:0] R3956;
  wire [63:0] R3955;
  wire [63:0] R3954;
  wire [31:0] R3953;
  wire [63:0] R3952;
  wire [63:0] R3951;
  wire [63:0] R3950;
  wire [63:0] R3949;
  wire [63:0] R3948;
  wire [63:0] R3947;
  wire [63:0] R3946;
  wire [31:0] R3945;
  wire [31:0] R3944;
  wire [31:0] R3943;
  wire [63:0] R3942;
  wire [63:0] R3941;
  wire [63:0] R3940;
  wire [63:0] R3939;
  wire [63:0] R3938;
  wire [63:0] R3937;
  wire [63:0] R3936;
  wire [63:0] R3935;
  wire [63:0] R3934;
  wire [63:0] R3933;
  wire [63:0] R3932;
  wire [63:0] R3931;
  wire [63:0] R3930;
  wire [63:0] R3929;
  wire [63:0] R3928;
  wire [63:0] R3927;
  wire [63:0] R3926;
  wire [63:0] R3925;
  wire [63:0] R3924;
  wire [63:0] R3923;
  wire [63:0] R3922;
  wire [63:0] R3921;
  wire [63:0] R3920;
  wire [63:0] R3919;
  wire [0:0] R3918;
  wire [0:0] R3917;
  wire [0:0] R3916;
  wire [0:0] R3915;
  wire [0:0] R3914;
  wire [0:0] R3913;
  wire [0:0] R3912;
  wire [0:0] R3911;
  wire [0:0] R3910;
  wire [0:0] R3909;
  wire [0:0] R3908;
  wire [0:0] R3907;
  wire [0:0] R3906;
  wire [0:0] R3905;
  wire [0:0] R3904;
  wire [0:0] R3903;
  wire [0:0] R3902;
  wire [0:0] R3901;
  wire [0:0] R3900;
  wire [0:0] R3899;
  wire [0:0] R3898;
  wire [0:0] R3897;
  wire [0:0] R3896;
  wire [0:0] R3895;
  wire [0:0] R3894;
  wire [0:0] R3893;
  wire [0:0] R3892;
  wire [0:0] R3891;
  wire [0:0] R3890;
  wire [0:0] R3889;
  wire [0:0] R3888;
  wire [0:0] R3887;
  wire [0:0] R3886;
  wire [0:0] R3885;
  wire [0:0] R3884;
  wire [0:0] R3883;
  wire [0:0] R3882;
  wire [0:0] R3881;
  wire [0:0] R3880;
  wire [0:0] R3879;
  wire [0:0] R3878;
  wire [0:0] R3877;
  wire [0:0] R3876;
  wire [0:0] R3875;
  wire [0:0] R3874;
  wire [0:0] R3873;
  wire [0:0] R3872;
  wire [0:0] R3871;
  wire [0:0] R3870;
  wire [0:0] R3869;
  wire [0:0] R3868;
  wire [0:0] R3867;
  wire [0:0] R3866;
  wire [0:0] R3865;
  wire [0:0] R3864;
  wire [0:0] R3863;
  wire [0:0] R3862;
  wire [0:0] R3861;
  wire [0:0] R3860;
  wire [0:0] R3859;
  wire [0:0] R3858;
  wire [0:0] R3857;
  wire [0:0] R3856;
  wire [0:0] R3855;
  wire [0:0] R3854;
  wire [0:0] R3853;
  wire [0:0] R3852;
  wire [0:0] R3851;
  wire [0:0] R3850;
  wire [0:0] R3849;
  wire [0:0] R3848;
  wire [0:0] R3847;
  wire [0:0] R3846;
  wire [0:0] R3845;
  wire [0:0] R3844;
  wire [0:0] R3843;
  wire [0:0] R3842;
  wire [0:0] R3841;
  wire [0:0] R3840;
  wire [0:0] R3839;
  wire [0:0] R3838;
  wire [0:0] R3837;
  wire [0:0] R3836;
  wire [0:0] R3835;
  wire [0:0] R3834;
  wire [0:0] R3833;
  wire [0:0] R3832;
  wire [0:0] R3831;
  wire [0:0] R3830;
  wire [0:0] R3829;
  wire [0:0] R3828;
  wire [0:0] R3827;
  wire [0:0] R3826;
  wire [0:0] R3825;
  wire [0:0] R3824;
  wire [0:0] R3823;
  wire [0:0] R3822;
  wire [0:0] R3821;
  wire [0:0] R3820;
  wire [0:0] R3819;
  wire [0:0] R3818;
  wire [0:0] R3817;
  wire [0:0] R3816;
  wire [0:0] R3815;
  wire [0:0] R3814;
  wire [0:0] R3813;
  wire [0:0] R3812;
  wire [0:0] R3811;
  wire [0:0] R3810;
  wire [0:0] R3809;
  wire [0:0] R3808;
  wire [0:0] R3807;
  wire [0:0] R3806;
  wire [0:0] R3805;
  wire [0:0] R3804;
  wire [0:0] R3803;
  wire [0:0] R3802;
  wire [0:0] R3801;
  wire [0:0] R3800;
  wire [0:0] R3799;
  wire [0:0] R3798;
  wire [0:0] R3797;
  wire [0:0] R3796;
  wire [0:0] R3795;
  wire [0:0] R3794;
  wire [0:0] R3793;
  wire [0:0] R3792;
  wire [0:0] R3791;
  wire [0:0] R3790;
  wire [0:0] R3789;
  wire [0:0] R3788;
  wire [0:0] R3787;
  wire [0:0] R3786;
  wire [0:0] R3785;
  wire [0:0] R3784;
  wire [0:0] R3783;
  wire [0:0] R3782;
  wire [0:0] R3781;
  wire [0:0] R3780;
  wire [0:0] R3779;
  wire [0:0] R3778;
  wire [0:0] R3777;
  wire [0:0] R3776;
  wire [0:0] R3775;
  wire [0:0] R3774;
  wire [0:0] R3773;
  wire [0:0] R3772;
  wire [0:0] R3771;
  wire [0:0] R3770;
  wire [0:0] R3769;
  wire [0:0] R3768;
  wire [0:0] R3767;
  wire [0:0] R3766;
  wire [0:0] R3765;
  wire [0:0] R3764;
  wire [0:0] R3763;
  wire [0:0] R3762;
  wire [0:0] R3761;
  wire [0:0] R3760;
  wire [0:0] R3759;
  wire [0:0] R3758;
  wire [0:0] R3757;
  wire [0:0] R3756;
  wire [0:0] R3755;
  wire [0:0] R3754;
  wire [0:0] R3753;
  wire [0:0] R3752;
  wire [0:0] R3751;
  wire [0:0] R3750;
  wire [0:0] R3749;
  wire [0:0] R3748;
  wire [0:0] R3747;
  wire [0:0] R3746;
  wire [0:0] R3745;
  wire [0:0] R3744;
  wire [0:0] R3743;
  wire [0:0] R3742;
  wire [0:0] R3741;
  wire [0:0] R3740;
  wire [0:0] R3739;
  wire [0:0] R3738;
  wire [0:0] R3737;
  wire [0:0] R3736;
  wire [0:0] R3735;
  wire [0:0] R3734;
  wire [0:0] R3733;
  wire [0:0] R3732;
  wire [0:0] R3731;
  wire [0:0] R3730;
  wire [0:0] R3729;
  wire [0:0] R3728;
  wire [0:0] R3727;
  wire [0:0] R3726;
  wire [0:0] R3725;
  wire [63:0] R3724;
  wire [31:0] R3723;
  wire [31:0] R3722;
  wire [31:0] R3721;
  wire [31:0] R3720;
  wire [31:0] R3719;
  wire [31:0] R3718;
  wire [31:0] R3717;
  wire [31:0] R3716;
  wire [31:0] R3715;
  wire [31:0] R3714;
  wire [31:0] R3713;
  wire [31:0] R3712;
  wire [31:0] R3711;
  wire [31:0] R3710;
  wire [31:0] R3709;
  wire [31:0] R3708;
  wire [31:0] R3707;
  wire [31:0] R3706;
  wire [31:0] R3705;
  wire [31:0] R3704;
  wire [31:0] R3703;
  wire [31:0] R3702;
  wire [31:0] R3701;
  wire [31:0] R3700;
  wire [31:0] R3699;
  wire [31:0] R3698;
  wire [31:0] R3697;
  wire [31:0] R3696;
  wire [31:0] R3695;
  wire [31:0] R3694;
  wire [31:0] R3693;
  wire [31:0] R3692;
  wire [31:0] R3691;
  wire [31:0] R3690;
  wire [31:0] R3689;
  wire [31:0] R3688;
  wire [31:0] R3687;
  wire [31:0] R3686;
  wire [31:0] R3685;
  wire [31:0] R3684;
  wire [31:0] R3683;
  wire [31:0] R3682;
  wire [31:0] R3681;
  wire [31:0] R3680;
  wire [31:0] R3679;
  wire [31:0] R3678;
  wire [31:0] R3677;
  wire [31:0] R3676;
  wire [31:0] R3675;
  wire [31:0] R3674;
  wire [31:0] R3673;
  wire [31:0] R3672;
  wire [31:0] R3671;
  wire [31:0] R3670;
  wire [31:0] R3669;
  wire [31:0] R3668;
  wire [31:0] R3667;
  wire [31:0] R3666;
  wire [31:0] R3665;
  wire [31:0] R3664;
  wire [31:0] R3663;
  wire [31:0] R3662;
  wire [31:0] R3661;
  wire [31:0] R3660;
  wire [31:0] R3659;
  wire [31:0] R3658;
  wire [31:0] R3657;
  wire [31:0] R3656;
  wire [31:0] R3655;
  wire [31:0] R3654;
  wire [31:0] R3653;
  wire [31:0] R3652;
  wire [31:0] R3651;
  wire [31:0] R3650;
  wire [31:0] R3649;
  wire [31:0] R3648;
  wire [31:0] R3647;
  wire [31:0] R3646;
  wire [31:0] R3645;
  wire [31:0] R3644;
  wire [31:0] R3643;
  wire [31:0] R3642;
  wire [31:0] R3641;
  wire [31:0] R3640;
  wire [31:0] R3639;
  wire [31:0] R3638;
  wire [31:0] R3637;
  wire [31:0] R3636;
  wire [31:0] R3635;
  wire [31:0] R3634;
  wire [31:0] R3633;
  wire [31:0] R3632;
  wire [31:0] R3631;
  wire [31:0] R3630;
  wire [31:0] R3629;
  wire [31:0] R3628;
  wire [31:0] R3627;
  wire [31:0] R3626;
  wire [31:0] R3625;
  wire [31:0] R3624;
  wire [31:0] R3623;
  wire [31:0] R3622;
  wire [31:0] R3621;
  wire [31:0] R3620;
  wire [31:0] R3619;
  wire [31:0] R3618;
  wire [31:0] R3617;
  wire [31:0] R3616;
  wire [31:0] R3615;
  wire [31:0] R3614;
  wire [31:0] R3613;
  wire [31:0] R3612;
  wire [31:0] R3611;
  wire [31:0] R3610;
  wire [31:0] R3609;
  wire [31:0] R3608;
  wire [31:0] R3607;
  wire [31:0] R3606;
  wire [31:0] R3605;
  wire [31:0] R3604;
  wire [31:0] R3603;
  wire [31:0] R3602;
  wire [31:0] R3601;
  wire [31:0] R3600;
  wire [31:0] R3599;
  wire [31:0] R3598;
  wire [31:0] R3597;
  wire [31:0] R3596;
  wire [31:0] R3595;
  wire [31:0] R3594;
  wire [31:0] R3593;
  wire [31:0] R3592;
  wire [31:0] R3591;
  wire [31:0] R3590;
  wire [31:0] R3589;
  wire [31:0] R3588;
  wire [31:0] R3587;
  wire [31:0] R3586;
  wire [31:0] R3585;
  wire [31:0] R3584;
  wire [31:0] R3583;
  wire [31:0] R3582;
  wire [31:0] R3581;
  wire [31:0] R3580;
  wire [31:0] R3579;
  wire [31:0] R3578;
  wire [31:0] R3577;
  wire [31:0] R3576;
  wire [31:0] R3575;
  wire [31:0] R3574;
  wire [31:0] R3573;
  wire [31:0] R3572;
  wire [31:0] R3571;
  wire [31:0] R3570;
  wire [31:0] R3569;
  wire [31:0] R3568;
  wire [31:0] R3567;
  wire [31:0] R3566;
  wire [31:0] R3565;
  wire [31:0] R3564;
  wire [31:0] R3563;
  wire [31:0] R3562;
  wire [31:0] R3561;
  wire [31:0] R3560;
  wire [31:0] R3559;
  wire [31:0] R3558;
  wire [31:0] R3557;
  wire [31:0] R3556;
  wire [31:0] R3555;
  wire [31:0] R3554;
  wire [31:0] R3553;
  wire [31:0] R3552;
  wire [31:0] R3551;
  wire [31:0] R3550;
  wire [31:0] R3549;
  wire [31:0] R3548;
  wire [31:0] R3547;
  wire [31:0] R3546;
  wire [31:0] R3545;
  wire [31:0] R3544;
  wire [31:0] R3543;
  wire [31:0] R3542;
  wire [31:0] R3541;
  wire [31:0] R3540;
  wire [31:0] R3539;
  wire [31:0] R3538;
  wire [31:0] R3537;
  wire [31:0] R3536;
  wire [63:0] R3535;
  wire [63:0] R3534;
  wire [63:0] R3533;
  wire [31:0] R3532;
  wire [31:0] R3531;
  wire [31:0] R3530;
  wire [31:0] R3529;
  wire [31:0] R3528;
  wire [31:0] R3527;
  wire [31:0] R3526;
  wire [31:0] R3525;
  wire [31:0] R3524;
  wire [31:0] R3523;
  wire [31:0] R3522;
  wire [31:0] R3521;
  wire [31:0] R3520;
  wire [31:0] R3519;
  wire [31:0] R3518;
  wire [31:0] R3517;
  wire [31:0] R3516;
  wire [31:0] R3515;
  wire [31:0] R3514;
  wire [31:0] R3513;
  wire [31:0] R3512;
  wire [31:0] R3511;
  wire [31:0] R3510;
  wire [31:0] R3509;
  wire [31:0] R3508;
  wire [31:0] R3507;
  wire [31:0] R3506;
  wire [31:0] R3505;
  wire [31:0] R3504;
  wire [31:0] R3503;
  wire [31:0] R3502;
  wire [31:0] R3501;
  wire [31:0] R3500;
  wire [31:0] R3499;
  wire [31:0] R3498;
  wire [31:0] R3497;
  wire [31:0] R3496;
  wire [31:0] R3495;
  wire [31:0] R3494;
  wire [31:0] R3493;
  wire [31:0] R3492;
  wire [31:0] R3491;
  wire [31:0] R3490;
  wire [31:0] R3489;
  wire [31:0] R3488;
  wire [31:0] R3487;
  wire [31:0] R3486;
  wire [31:0] R3485;
  wire [31:0] R3484;
  wire [31:0] R3483;
  wire [31:0] R3482;
  wire [31:0] R3481;
  wire [31:0] R3480;
  wire [31:0] R3479;
  wire [31:0] R3478;
  wire [31:0] R3477;
  wire [31:0] R3476;
  wire [31:0] R3475;
  wire [31:0] R3474;
  wire [31:0] R3473;
  wire [31:0] R3472;
  wire [31:0] R3471;
  wire [31:0] R3470;
  wire [31:0] R3469;
  wire [31:0] R3468;
  wire [31:0] R3467;
  wire [31:0] R3466;
  wire [31:0] R3465;
  wire [31:0] R3464;
  wire [31:0] R3463;
  wire [31:0] R3462;
  wire [31:0] R3461;
  wire [31:0] R3460;
  wire [31:0] R3459;
  wire [31:0] R3458;
  wire [31:0] R3457;
  wire [31:0] R3456;
  wire [31:0] R3455;
  wire [31:0] R3454;
  wire [31:0] R3453;
  wire [31:0] R3452;
  wire [31:0] R3451;
  wire [31:0] R3450;
  wire [31:0] R3449;
  wire [31:0] R3448;
  wire [31:0] R3447;
  wire [31:0] R3446;
  wire [31:0] R3445;
  wire [31:0] R3444;
  wire [31:0] R3443;
  wire [31:0] R3442;
  wire [31:0] R3441;
  wire [31:0] R3440;
  wire [31:0] R3439;
  wire [31:0] R3438;
  wire [31:0] R3437;
  wire [31:0] R3436;
  wire [31:0] R3435;
  wire [31:0] R3434;
  wire [31:0] R3433;
  wire [31:0] R3432;
  wire [31:0] R3431;
  wire [31:0] R3430;
  wire [31:0] R3429;
  wire [31:0] R3428;
  wire [31:0] R3427;
  wire [31:0] R3426;
  wire [31:0] R3425;
  wire [31:0] R3424;
  wire [31:0] R3423;
  wire [31:0] R3422;
  wire [31:0] R3421;
  wire [31:0] R3420;
  wire [31:0] R3419;
  wire [31:0] R3418;
  wire [31:0] R3417;
  wire [31:0] R3416;
  wire [31:0] R3415;
  wire [31:0] R3414;
  wire [31:0] R3413;
  wire [31:0] R3412;
  wire [31:0] R3411;
  wire [31:0] R3410;
  wire [31:0] R3409;
  wire [31:0] R3408;
  wire [31:0] R3407;
  wire [31:0] R3406;
  wire [31:0] R3405;
  wire [31:0] R3404;
  wire [31:0] R3403;
  wire [31:0] R3402;
  wire [31:0] R3401;
  wire [31:0] R3400;
  wire [31:0] R3399;
  wire [31:0] R3398;
  wire [31:0] R3397;
  wire [31:0] R3396;
  wire [31:0] R3395;
  wire [31:0] R3394;
  wire [31:0] R3393;
  wire [31:0] R3392;
  wire [31:0] R3391;
  wire [31:0] R3390;
  wire [31:0] R3389;
  wire [31:0] R3388;
  wire [31:0] R3387;
  wire [31:0] R3386;
  wire [31:0] R3385;
  wire [31:0] R3384;
  wire [31:0] R3383;
  wire [31:0] R3382;
  wire [31:0] R3381;
  wire [31:0] R3380;
  wire [31:0] R3379;
  wire [31:0] R3378;
  wire [31:0] R3377;
  wire [31:0] R3376;
  wire [31:0] R3375;
  wire [31:0] R3374;
  wire [31:0] R3373;
  wire [31:0] R3372;
  wire [31:0] R3371;
  wire [31:0] R3370;
  wire [31:0] R3369;
  wire [31:0] R3368;
  wire [31:0] R3367;
  wire [31:0] R3366;
  wire [31:0] R3365;
  wire [31:0] R3364;
  wire [31:0] R3363;
  wire [31:0] R3362;
  wire [31:0] R3361;
  wire [31:0] R3360;
  wire [31:0] R3359;
  wire [31:0] R3358;
  wire [31:0] R3357;
  wire [31:0] R3356;
  wire [31:0] R3355;
  wire [31:0] R3354;
  wire [31:0] R3353;
  wire [31:0] R3352;
  wire [31:0] R3351;
  wire [31:0] R3350;
  wire [31:0] R3349;
  wire [31:0] R3348;
  wire [31:0] R3347;
  wire [31:0] R3346;
  wire [31:0] R3345;
  wire [31:0] R3344;
  wire [31:0] R3343;
  wire [31:0] R3342;
  wire [31:0] R3341;
  wire [31:0] R3340;
  wire [31:0] R3339;
  wire [31:0] R3338;
  wire [63:0] R3337;
  wire [31:0] R3336;
  wire [31:0] R3335;
  wire [63:0] R3334;
  wire [31:0] R3333;
  wire [63:0] R3332;
  wire [63:0] R3331;
  wire [63:0] R3330;
  wire [63:0] R3329;
  wire [63:0] R3328;
  wire [63:0] R3327;
  wire [31:0] R3326;
  wire [63:0] R3325;
  wire [63:0] R3324;
  wire [63:0] R3323;
  wire [63:0] R3322;
  wire [63:0] R3321;
  wire [63:0] R3320;
  wire [63:0] R3319;
  wire [31:0] R3318;
  wire [31:0] R3317;
  wire [31:0] R3316;
  wire [63:0] R3315;
  wire [63:0] R3314;
  wire [63:0] R3313;
  wire [63:0] R3312;
  wire [63:0] R3311;
  wire [63:0] R3310;
  wire [63:0] R3309;
  wire [63:0] R3308;
  wire [63:0] R3307;
  wire [63:0] R3306;
  wire [63:0] R3305;
  wire [63:0] R3304;
  wire [63:0] R3303;
  wire [63:0] R3302;
  wire [63:0] R3301;
  wire [63:0] R3300;
  wire [63:0] R3299;
  wire [63:0] R3298;
  wire [63:0] R3297;
  wire [63:0] R3296;
  wire [63:0] R3295;
  wire [63:0] R3294;
  wire [63:0] R3293;
  wire [63:0] R3292;
  wire [0:0] R3291;
  wire [0:0] R3290;
  wire [0:0] R3289;
  wire [0:0] R3288;
  wire [0:0] R3287;
  wire [0:0] R3286;
  wire [0:0] R3285;
  wire [0:0] R3284;
  wire [0:0] R3283;
  wire [0:0] R3282;
  wire [0:0] R3281;
  wire [0:0] R3280;
  wire [0:0] R3279;
  wire [0:0] R3278;
  wire [0:0] R3277;
  wire [0:0] R3276;
  wire [0:0] R3275;
  wire [0:0] R3274;
  wire [0:0] R3273;
  wire [0:0] R3272;
  wire [0:0] R3271;
  wire [0:0] R3270;
  wire [0:0] R3269;
  wire [0:0] R3268;
  wire [0:0] R3267;
  wire [0:0] R3266;
  wire [0:0] R3265;
  wire [0:0] R3264;
  wire [0:0] R3263;
  wire [0:0] R3262;
  wire [0:0] R3261;
  wire [0:0] R3260;
  wire [0:0] R3259;
  wire [0:0] R3258;
  wire [0:0] R3257;
  wire [0:0] R3256;
  wire [0:0] R3255;
  wire [0:0] R3254;
  wire [0:0] R3253;
  wire [0:0] R3252;
  wire [0:0] R3251;
  wire [0:0] R3250;
  wire [0:0] R3249;
  wire [0:0] R3248;
  wire [0:0] R3247;
  wire [0:0] R3246;
  wire [0:0] R3245;
  wire [0:0] R3244;
  wire [0:0] R3243;
  wire [0:0] R3242;
  wire [0:0] R3241;
  wire [0:0] R3240;
  wire [0:0] R3239;
  wire [0:0] R3238;
  wire [0:0] R3237;
  wire [0:0] R3236;
  wire [0:0] R3235;
  wire [0:0] R3234;
  wire [0:0] R3233;
  wire [0:0] R3232;
  wire [0:0] R3231;
  wire [0:0] R3230;
  wire [0:0] R3229;
  wire [0:0] R3228;
  wire [0:0] R3227;
  wire [0:0] R3226;
  wire [0:0] R3225;
  wire [0:0] R3224;
  wire [0:0] R3223;
  wire [0:0] R3222;
  wire [0:0] R3221;
  wire [0:0] R3220;
  wire [0:0] R3219;
  wire [0:0] R3218;
  wire [0:0] R3217;
  wire [0:0] R3216;
  wire [0:0] R3215;
  wire [0:0] R3214;
  wire [0:0] R3213;
  wire [0:0] R3212;
  wire [0:0] R3211;
  wire [0:0] R3210;
  wire [0:0] R3209;
  wire [0:0] R3208;
  wire [0:0] R3207;
  wire [0:0] R3206;
  wire [0:0] R3205;
  wire [0:0] R3204;
  wire [0:0] R3203;
  wire [0:0] R3202;
  wire [0:0] R3201;
  wire [0:0] R3200;
  wire [0:0] R3199;
  wire [0:0] R3198;
  wire [0:0] R3197;
  wire [0:0] R3196;
  wire [0:0] R3195;
  wire [0:0] R3194;
  wire [0:0] R3193;
  wire [0:0] R3192;
  wire [0:0] R3191;
  wire [0:0] R3190;
  wire [0:0] R3189;
  wire [0:0] R3188;
  wire [0:0] R3187;
  wire [0:0] R3186;
  wire [0:0] R3185;
  wire [0:0] R3184;
  wire [0:0] R3183;
  wire [0:0] R3182;
  wire [0:0] R3181;
  wire [0:0] R3180;
  wire [0:0] R3179;
  wire [0:0] R3178;
  wire [0:0] R3177;
  wire [0:0] R3176;
  wire [0:0] R3175;
  wire [0:0] R3174;
  wire [0:0] R3173;
  wire [0:0] R3172;
  wire [0:0] R3171;
  wire [0:0] R3170;
  wire [0:0] R3169;
  wire [0:0] R3168;
  wire [0:0] R3167;
  wire [0:0] R3166;
  wire [0:0] R3165;
  wire [0:0] R3164;
  wire [0:0] R3163;
  wire [0:0] R3162;
  wire [0:0] R3161;
  wire [0:0] R3160;
  wire [0:0] R3159;
  wire [0:0] R3158;
  wire [0:0] R3157;
  wire [0:0] R3156;
  wire [0:0] R3155;
  wire [0:0] R3154;
  wire [0:0] R3153;
  wire [0:0] R3152;
  wire [0:0] R3151;
  wire [0:0] R3150;
  wire [0:0] R3149;
  wire [0:0] R3148;
  wire [0:0] R3147;
  wire [0:0] R3146;
  wire [0:0] R3145;
  wire [0:0] R3144;
  wire [0:0] R3143;
  wire [0:0] R3142;
  wire [0:0] R3141;
  wire [0:0] R3140;
  wire [0:0] R3139;
  wire [0:0] R3138;
  wire [0:0] R3137;
  wire [0:0] R3136;
  wire [0:0] R3135;
  wire [0:0] R3134;
  wire [0:0] R3133;
  wire [0:0] R3132;
  wire [0:0] R3131;
  wire [0:0] R3130;
  wire [0:0] R3129;
  wire [0:0] R3128;
  wire [0:0] R3127;
  wire [0:0] R3126;
  wire [0:0] R3125;
  wire [0:0] R3124;
  wire [0:0] R3123;
  wire [0:0] R3122;
  wire [0:0] R3121;
  wire [0:0] R3120;
  wire [0:0] R3119;
  wire [0:0] R3118;
  wire [0:0] R3117;
  wire [0:0] R3116;
  wire [0:0] R3115;
  wire [0:0] R3114;
  wire [0:0] R3113;
  wire [0:0] R3112;
  wire [0:0] R3111;
  wire [0:0] R3110;
  wire [0:0] R3109;
  wire [0:0] R3108;
  wire [0:0] R3107;
  wire [0:0] R3106;
  wire [0:0] R3105;
  wire [0:0] R3104;
  wire [0:0] R3103;
  wire [0:0] R3102;
  wire [0:0] R3101;
  wire [0:0] R3100;
  wire [0:0] R3099;
  wire [0:0] R3098;
  wire [0:0] R3097;
  wire [0:0] R3096;
  wire [0:0] R3095;
  wire [0:0] R3094;
  wire [0:0] R3093;
  wire [0:0] R3092;
  wire [0:0] R3091;
  wire [0:0] R3090;
  wire [0:0] R3089;
  wire [0:0] R3088;
  wire [0:0] R3087;
  wire [0:0] R3086;
  wire [0:0] R3085;
  wire [0:0] R3084;
  wire [63:0] R3083;
  wire [31:0] R3082;
  wire [31:0] R3081;
  wire [31:0] R3080;
  wire [31:0] R3079;
  wire [31:0] R3078;
  wire [31:0] R3077;
  wire [31:0] R3076;
  wire [31:0] R3075;
  wire [31:0] R3074;
  wire [31:0] R3073;
  wire [31:0] R3072;
  wire [31:0] R3071;
  wire [31:0] R3070;
  wire [31:0] R3069;
  wire [31:0] R3068;
  wire [31:0] R3067;
  wire [31:0] R3066;
  wire [31:0] R3065;
  wire [31:0] R3064;
  wire [31:0] R3063;
  wire [31:0] R3062;
  wire [31:0] R3061;
  wire [31:0] R3060;
  wire [31:0] R3059;
  wire [31:0] R3058;
  wire [31:0] R3057;
  wire [31:0] R3056;
  wire [31:0] R3055;
  wire [31:0] R3054;
  wire [31:0] R3053;
  wire [31:0] R3052;
  wire [31:0] R3051;
  wire [31:0] R3050;
  wire [31:0] R3049;
  wire [31:0] R3048;
  wire [31:0] R3047;
  wire [31:0] R3046;
  wire [31:0] R3045;
  wire [31:0] R3044;
  wire [31:0] R3043;
  wire [31:0] R3042;
  wire [31:0] R3041;
  wire [31:0] R3040;
  wire [31:0] R3039;
  wire [31:0] R3038;
  wire [31:0] R3037;
  wire [31:0] R3036;
  wire [31:0] R3035;
  wire [31:0] R3034;
  wire [31:0] R3033;
  wire [31:0] R3032;
  wire [31:0] R3031;
  wire [31:0] R3030;
  wire [31:0] R3029;
  wire [31:0] R3028;
  wire [31:0] R3027;
  wire [31:0] R3026;
  wire [31:0] R3025;
  wire [31:0] R3024;
  wire [31:0] R3023;
  wire [31:0] R3022;
  wire [31:0] R3021;
  wire [31:0] R3020;
  wire [31:0] R3019;
  wire [31:0] R3018;
  wire [31:0] R3017;
  wire [31:0] R3016;
  wire [31:0] R3015;
  wire [31:0] R3014;
  wire [31:0] R3013;
  wire [31:0] R3012;
  wire [31:0] R3011;
  wire [31:0] R3010;
  wire [31:0] R3009;
  wire [31:0] R3008;
  wire [31:0] R3007;
  wire [31:0] R3006;
  wire [31:0] R3005;
  wire [31:0] R3004;
  wire [31:0] R3003;
  wire [31:0] R3002;
  wire [31:0] R3001;
  wire [31:0] R3000;
  wire [31:0] R2999;
  wire [31:0] R2998;
  wire [31:0] R2997;
  wire [31:0] R2996;
  wire [31:0] R2995;
  wire [31:0] R2994;
  wire [31:0] R2993;
  wire [31:0] R2992;
  wire [31:0] R2991;
  wire [31:0] R2990;
  wire [31:0] R2989;
  wire [31:0] R2988;
  wire [31:0] R2987;
  wire [31:0] R2986;
  wire [31:0] R2985;
  wire [31:0] R2984;
  wire [31:0] R2983;
  wire [31:0] R2982;
  wire [31:0] R2981;
  wire [31:0] R2980;
  wire [31:0] R2979;
  wire [31:0] R2978;
  wire [31:0] R2977;
  wire [31:0] R2976;
  wire [31:0] R2975;
  wire [31:0] R2974;
  wire [31:0] R2973;
  wire [31:0] R2972;
  wire [31:0] R2971;
  wire [31:0] R2970;
  wire [31:0] R2969;
  wire [31:0] R2968;
  wire [31:0] R2967;
  wire [31:0] R2966;
  wire [31:0] R2965;
  wire [31:0] R2964;
  wire [31:0] R2963;
  wire [31:0] R2962;
  wire [31:0] R2961;
  wire [31:0] R2960;
  wire [31:0] R2959;
  wire [31:0] R2958;
  wire [31:0] R2957;
  wire [31:0] R2956;
  wire [31:0] R2955;
  wire [31:0] R2954;
  wire [31:0] R2953;
  wire [31:0] R2952;
  wire [31:0] R2951;
  wire [31:0] R2950;
  wire [31:0] R2949;
  wire [31:0] R2948;
  wire [31:0] R2947;
  wire [31:0] R2946;
  wire [31:0] R2945;
  wire [31:0] R2944;
  wire [31:0] R2943;
  wire [31:0] R2942;
  wire [31:0] R2941;
  wire [31:0] R2940;
  wire [31:0] R2939;
  wire [31:0] R2938;
  wire [31:0] R2937;
  wire [31:0] R2936;
  wire [31:0] R2935;
  wire [31:0] R2934;
  wire [31:0] R2933;
  wire [31:0] R2932;
  wire [31:0] R2931;
  wire [31:0] R2930;
  wire [31:0] R2929;
  wire [31:0] R2928;
  wire [31:0] R2927;
  wire [31:0] R2926;
  wire [31:0] R2925;
  wire [31:0] R2924;
  wire [31:0] R2923;
  wire [31:0] R2922;
  wire [31:0] R2921;
  wire [31:0] R2920;
  wire [31:0] R2919;
  wire [31:0] R2918;
  wire [31:0] R2917;
  wire [31:0] R2916;
  wire [31:0] R2915;
  wire [31:0] R2914;
  wire [31:0] R2913;
  wire [31:0] R2912;
  wire [31:0] R2911;
  wire [31:0] R2910;
  wire [31:0] R2909;
  wire [31:0] R2908;
  wire [31:0] R2907;
  wire [31:0] R2906;
  wire [31:0] R2905;
  wire [31:0] R2904;
  wire [31:0] R2903;
  wire [31:0] R2902;
  wire [31:0] R2901;
  wire [31:0] R2900;
  wire [31:0] R2899;
  wire [31:0] R2898;
  wire [31:0] R2897;
  wire [31:0] R2896;
  wire [31:0] R2895;
  wire [31:0] R2894;
  wire [31:0] R2893;
  wire [31:0] R2892;
  wire [31:0] R2891;
  wire [31:0] R2890;
  wire [31:0] R2889;
  wire [31:0] R2888;
  wire [31:0] R2887;
  wire [31:0] R2886;
  wire [31:0] R2885;
  wire [31:0] R2884;
  wire [31:0] R2883;
  wire [31:0] R2882;
  wire [31:0] R2881;
  wire [63:0] R2880;
  wire [63:0] R2879;
  wire [63:0] R2878;
  wire [31:0] R2877;
  wire [31:0] R2876;
  wire [31:0] R2875;
  wire [31:0] R2874;
  wire [31:0] R2873;
  wire [31:0] R2872;
  wire [31:0] R2871;
  wire [31:0] R2870;
  wire [31:0] R2869;
  wire [31:0] R2868;
  wire [31:0] R2867;
  wire [31:0] R2866;
  wire [31:0] R2865;
  wire [31:0] R2864;
  wire [31:0] R2863;
  wire [31:0] R2862;
  wire [31:0] R2861;
  wire [31:0] R2860;
  wire [31:0] R2859;
  wire [31:0] R2858;
  wire [31:0] R2857;
  wire [31:0] R2856;
  wire [31:0] R2855;
  wire [31:0] R2854;
  wire [31:0] R2853;
  wire [31:0] R2852;
  wire [31:0] R2851;
  wire [31:0] R2850;
  wire [31:0] R2849;
  wire [31:0] R2848;
  wire [31:0] R2847;
  wire [31:0] R2846;
  wire [31:0] R2845;
  wire [31:0] R2844;
  wire [31:0] R2843;
  wire [31:0] R2842;
  wire [31:0] R2841;
  wire [31:0] R2840;
  wire [31:0] R2839;
  wire [31:0] R2838;
  wire [31:0] R2837;
  wire [31:0] R2836;
  wire [31:0] R2835;
  wire [31:0] R2834;
  wire [31:0] R2833;
  wire [31:0] R2832;
  wire [31:0] R2831;
  wire [31:0] R2830;
  wire [31:0] R2829;
  wire [31:0] R2828;
  wire [31:0] R2827;
  wire [31:0] R2826;
  wire [31:0] R2825;
  wire [31:0] R2824;
  wire [31:0] R2823;
  wire [31:0] R2822;
  wire [31:0] R2821;
  wire [31:0] R2820;
  wire [31:0] R2819;
  wire [31:0] R2818;
  wire [31:0] R2817;
  wire [31:0] R2816;
  wire [31:0] R2815;
  wire [31:0] R2814;
  wire [31:0] R2813;
  wire [31:0] R2812;
  wire [31:0] R2811;
  wire [31:0] R2810;
  wire [31:0] R2809;
  wire [31:0] R2808;
  wire [31:0] R2807;
  wire [31:0] R2806;
  wire [31:0] R2805;
  wire [31:0] R2804;
  wire [31:0] R2803;
  wire [31:0] R2802;
  wire [31:0] R2801;
  wire [31:0] R2800;
  wire [31:0] R2799;
  wire [31:0] R2798;
  wire [31:0] R2797;
  wire [31:0] R2796;
  wire [31:0] R2795;
  wire [31:0] R2794;
  wire [31:0] R2793;
  wire [31:0] R2792;
  wire [31:0] R2791;
  wire [31:0] R2790;
  wire [31:0] R2789;
  wire [31:0] R2788;
  wire [31:0] R2787;
  wire [31:0] R2786;
  wire [31:0] R2785;
  wire [31:0] R2784;
  wire [31:0] R2783;
  wire [31:0] R2782;
  wire [31:0] R2781;
  wire [31:0] R2780;
  wire [31:0] R2779;
  wire [31:0] R2778;
  wire [31:0] R2777;
  wire [31:0] R2776;
  wire [31:0] R2775;
  wire [31:0] R2774;
  wire [31:0] R2773;
  wire [31:0] R2772;
  wire [31:0] R2771;
  wire [31:0] R2770;
  wire [31:0] R2769;
  wire [31:0] R2768;
  wire [31:0] R2767;
  wire [31:0] R2766;
  wire [31:0] R2765;
  wire [31:0] R2764;
  wire [31:0] R2763;
  wire [31:0] R2762;
  wire [31:0] R2761;
  wire [31:0] R2760;
  wire [31:0] R2759;
  wire [31:0] R2758;
  wire [31:0] R2757;
  wire [31:0] R2756;
  wire [31:0] R2755;
  wire [31:0] R2754;
  wire [31:0] R2753;
  wire [31:0] R2752;
  wire [31:0] R2751;
  wire [31:0] R2750;
  wire [31:0] R2749;
  wire [31:0] R2748;
  wire [31:0] R2747;
  wire [31:0] R2746;
  wire [31:0] R2745;
  wire [31:0] R2744;
  wire [31:0] R2743;
  wire [31:0] R2742;
  wire [31:0] R2741;
  wire [31:0] R2740;
  wire [31:0] R2739;
  wire [31:0] R2738;
  wire [31:0] R2737;
  wire [31:0] R2736;
  wire [31:0] R2735;
  wire [31:0] R2734;
  wire [31:0] R2733;
  wire [31:0] R2732;
  wire [31:0] R2731;
  wire [31:0] R2730;
  wire [31:0] R2729;
  wire [31:0] R2728;
  wire [31:0] R2727;
  wire [31:0] R2726;
  wire [31:0] R2725;
  wire [31:0] R2724;
  wire [31:0] R2723;
  wire [31:0] R2722;
  wire [31:0] R2721;
  wire [31:0] R2720;
  wire [31:0] R2719;
  wire [31:0] R2718;
  wire [31:0] R2717;
  wire [31:0] R2716;
  wire [31:0] R2715;
  wire [31:0] R2714;
  wire [31:0] R2713;
  wire [31:0] R2712;
  wire [31:0] R2711;
  wire [31:0] R2710;
  wire [31:0] R2709;
  wire [31:0] R2708;
  wire [31:0] R2707;
  wire [31:0] R2706;
  wire [31:0] R2705;
  wire [31:0] R2704;
  wire [31:0] R2703;
  wire [31:0] R2702;
  wire [31:0] R2701;
  wire [31:0] R2700;
  wire [31:0] R2699;
  wire [31:0] R2698;
  wire [31:0] R2697;
  wire [31:0] R2696;
  wire [31:0] R2695;
  wire [31:0] R2694;
  wire [31:0] R2693;
  wire [31:0] R2692;
  wire [31:0] R2691;
  wire [31:0] R2690;
  wire [31:0] R2689;
  wire [31:0] R2688;
  wire [31:0] R2687;
  wire [31:0] R2686;
  wire [31:0] R2685;
  wire [31:0] R2684;
  wire [31:0] R2683;
  wire [31:0] R2682;
  wire [31:0] R2681;
  wire [31:0] R2680;
  wire [31:0] R2679;
  wire [31:0] R2678;
  wire [31:0] R2677;
  wire [31:0] R2676;
  wire [31:0] R2675;
  wire [31:0] R2674;
  wire [31:0] R2673;
  wire [31:0] R2672;
  wire [31:0] R2671;
  wire [31:0] R2670;
  wire [31:0] R2669;
  wire [7:0] mux28;
  wire [7:0] mux27;
  wire [7:0] mux26;
  wire [7:0] mux25;
  wire [7:0] mux24;
  wire [7:0] mux23;
  wire [7:0] mux22;
  wire [7:0] mux21;
  wire [7:0] mux20;
  wire [7:0] mux19;
  wire [7:0] mux18;
  wire [7:0] mux17;
  wire [7:0] mux16;
  wire [7:0] mux15;
  wire [7:0] mux14;
  wire [7:0] mux13;
  wire [7:0] mux12;
  wire [7:0] mux11;
  wire [7:0] mux10;
  wire [7:0] mux9;
  wire [7:0] mux8;
  wire [7:0] mux7;
  wire [7:0] mux6;
  wire [7:0] mux5;
  wire [7:0] mux4;
  wire [7:0] mux3;
  wire [7:0] mux2;
  wire [7:0] mux1;
  wire [7:0] mux0;
  wire [7:0] _2673;
  wire [7:0] _2532;
  wire [63:0] _2520;
  wire [63:0] _2519;
  wire [31:0] n_idx_2530;
  wire [31:0] _2518;
  wire [63:0] _2517;
  wire [63:0] _2516;
  wire [63:0] _2515;
  wire [63:0] _2514;
  wire [63:0] _2513;
  wire [63:0] _2512;
  wire [63:0] _2511;
  wire [63:0] _2510;
  wire [63:0] _2509;
  wire [63:0] _2508;
  wire [63:0] _2507;
  wire [63:0] _2506;
  wire [31:0] _2505;
  wire [63:0] _2504;
  wire [63:0] _2503;
  wire [63:0] _2502;
  wire [63:0] _2501;
  wire [63:0] _2500;
  wire [31:0] _2499;
  wire [63:0] _2498;
  wire [63:0] _2497;
  wire [63:0] _2496;
  wire [63:0] _2495;
  wire [63:0] _2494;
  wire [63:0] _2493;
  wire [63:0] _2492;
  wire [63:0] _2491;
  wire [63:0] _2490;
  wire [31:0] _2489;
  wire [63:0] _2488;
  wire [63:0] _2487;
  wire [63:0] _2486;
  wire [63:0] _2485;
  wire [63:0] _2484;
  wire [31:0] _2483;
  wire [63:0] _2482;
  wire [63:0] _2481;
  wire [63:0] _2480;
  wire [63:0] _2479;
  wire [63:0] _2478;
  wire [63:0] _2477;
  wire [63:0] _2476;
  wire [63:0] _2475;
  wire [63:0] _2474;
  wire [63:0] _2473;
  wire [63:0] _2472;
  wire [31:0] _2471;
  wire [63:0] _2470;
  wire [63:0] _2469;
  wire [63:0] _2468;
  wire [63:0] _2467;
  wire [63:0] _2466;
  wire [31:0] _2465;
  wire [63:0] _2464;
  wire [63:0] _2463;
  wire [63:0] _2462;
  wire [63:0] _2461;
  wire [63:0] _2460;
  wire [63:0] _2459;
  wire [63:0] _2458;
  wire [63:0] _2457;
  wire [63:0] _2456;
  wire [31:0] _2455;
  wire [63:0] _2454;
  wire [63:0] _2453;
  wire [63:0] _2452;
  wire [63:0] _2451;
  wire [63:0] _2450;
  wire [31:0] _2449;
  wire [63:0] _2448;
  wire [63:0] _2447;
  wire [63:0] _2446;
  wire [63:0] _2445;
  wire [31:0] _2444;
  wire [63:0] _2443;
  wire [63:0] _2442;
  wire [63:0] _2441;
  wire [0:0] ifout2555;
  wire [63:0] _2440;
  wire [63:0] _2439;
  wire [63:0] _2438;
  wire [63:0] _2437;
  wire [63:0] _2436;
  wire [63:0] _2435;
  wire [7:0] _2542;
  wire [63:0] _2434;
  wire [63:0] _2433;
  wire [31:0] n_idx_2541;
  wire [31:0] _2432;
  wire [63:0] _2431;
  wire [63:0] _2430;
  wire [63:0] _2429;
  wire [63:0] _2428;
  wire [63:0] _2427;
  wire [63:0] _2426;
  wire [63:0] _2425;
  wire [63:0] _2424;
  wire [63:0] _2423;
  wire [63:0] _2422;
  wire [63:0] _2421;
  wire [63:0] _2420;
  wire [31:0] _2419;
  wire [63:0] _2418;
  wire [63:0] _2417;
  wire [63:0] _2416;
  wire [63:0] _2415;
  wire [63:0] _2414;
  wire [31:0] _2413;
  wire [63:0] _2412;
  wire [63:0] _2411;
  wire [63:0] _2410;
  wire [63:0] _2409;
  wire [63:0] _2408;
  wire [63:0] _2407;
  wire [63:0] _2406;
  wire [63:0] _2405;
  wire [63:0] _2404;
  wire [31:0] _2403;
  wire [63:0] _2402;
  wire [63:0] _2401;
  wire [63:0] _2400;
  wire [63:0] _2399;
  wire [63:0] _2398;
  wire [31:0] _2397;
  wire [63:0] _2396;
  wire [63:0] _2395;
  wire [63:0] _2394;
  wire [63:0] _2393;
  wire [63:0] _2392;
  wire [63:0] _2391;
  wire [63:0] _2390;
  wire [63:0] _2389;
  wire [63:0] _2388;
  wire [63:0] _2387;
  wire [63:0] _2386;
  wire [31:0] _2385;
  wire [63:0] _2384;
  wire [63:0] _2383;
  wire [63:0] _2382;
  wire [63:0] _2381;
  wire [63:0] _2380;
  wire [31:0] _2379;
  wire [63:0] _2378;
  wire [63:0] _2377;
  wire [63:0] _2376;
  wire [63:0] _2375;
  wire [63:0] _2374;
  wire [63:0] _2373;
  wire [63:0] _2372;
  wire [63:0] _2371;
  wire [63:0] _2370;
  wire [31:0] _2369;
  wire [63:0] _2368;
  wire [63:0] _2367;
  wire [63:0] _2366;
  wire [63:0] _2365;
  wire [63:0] _2364;
  wire [31:0] _2363;
  wire [63:0] _2362;
  wire [63:0] _2361;
  wire [63:0] _2360;
  wire [63:0] _2359;
  wire [31:0] _2358;
  wire [63:0] _2357;
  wire [63:0] _2356;
  wire [63:0] _2355;
  wire [0:0] ifout2466;
  wire [63:0] _2354;
  wire [63:0] _2353;
  wire [63:0] _2352;
  wire [63:0] _2351;
  wire [63:0] _2350;
  wire [63:0] _2349;
  wire [7:0] _2552;
  wire [63:0] _2348;
  wire [63:0] _2347;
  wire [31:0] n_idx_2551;
  wire [31:0] _2346;
  wire [63:0] _2345;
  wire [63:0] _2344;
  wire [63:0] _2343;
  wire [63:0] _2342;
  wire [63:0] _2341;
  wire [63:0] _2340;
  wire [63:0] _2339;
  wire [63:0] _2338;
  wire [63:0] _2337;
  wire [63:0] _2336;
  wire [63:0] _2335;
  wire [63:0] _2334;
  wire [31:0] _2333;
  wire [63:0] _2332;
  wire [63:0] _2331;
  wire [63:0] _2330;
  wire [63:0] _2329;
  wire [63:0] _2328;
  wire [31:0] _2327;
  wire [63:0] _2326;
  wire [63:0] _2325;
  wire [63:0] _2324;
  wire [63:0] _2323;
  wire [63:0] _2322;
  wire [63:0] _2321;
  wire [63:0] _2320;
  wire [63:0] _2319;
  wire [63:0] _2318;
  wire [31:0] _2317;
  wire [63:0] _2316;
  wire [63:0] _2315;
  wire [63:0] _2314;
  wire [63:0] _2313;
  wire [63:0] _2312;
  wire [31:0] _2311;
  wire [63:0] _2310;
  wire [63:0] _2309;
  wire [63:0] _2308;
  wire [63:0] _2307;
  wire [63:0] _2306;
  wire [63:0] _2305;
  wire [63:0] _2304;
  wire [63:0] _2303;
  wire [63:0] _2302;
  wire [63:0] _2301;
  wire [63:0] _2300;
  wire [31:0] _2299;
  wire [63:0] _2298;
  wire [63:0] _2297;
  wire [63:0] _2296;
  wire [63:0] _2295;
  wire [63:0] _2294;
  wire [31:0] _2293;
  wire [63:0] _2292;
  wire [63:0] _2291;
  wire [63:0] _2290;
  wire [63:0] _2289;
  wire [63:0] _2288;
  wire [63:0] _2287;
  wire [63:0] _2286;
  wire [63:0] _2285;
  wire [63:0] _2284;
  wire [31:0] _2283;
  wire [63:0] _2282;
  wire [63:0] _2281;
  wire [63:0] _2280;
  wire [63:0] _2279;
  wire [63:0] _2278;
  wire [31:0] _2277;
  wire [63:0] _2276;
  wire [63:0] _2275;
  wire [63:0] _2274;
  wire [63:0] _2273;
  wire [31:0] _2272;
  wire [63:0] _2271;
  wire [63:0] _2270;
  wire [63:0] _2269;
  wire [0:0] ifout2377;
  wire [63:0] _2268;
  wire [63:0] _2267;
  wire [63:0] _2266;
  wire [63:0] _2265;
  wire [63:0] _2264;
  wire [63:0] _2263;
  wire [7:0] _2562;
  wire [63:0] _2262;
  wire [63:0] _2261;
  wire [31:0] n_idx_2561;
  wire [31:0] _2260;
  wire [63:0] _2259;
  wire [63:0] _2258;
  wire [63:0] _2257;
  wire [63:0] _2256;
  wire [63:0] _2255;
  wire [63:0] _2254;
  wire [63:0] _2253;
  wire [63:0] _2252;
  wire [63:0] _2251;
  wire [63:0] _2250;
  wire [63:0] _2249;
  wire [63:0] _2248;
  wire [31:0] _2247;
  wire [63:0] _2246;
  wire [63:0] _2245;
  wire [63:0] _2244;
  wire [63:0] _2243;
  wire [63:0] _2242;
  wire [31:0] _2241;
  wire [63:0] _2240;
  wire [63:0] _2239;
  wire [63:0] _2238;
  wire [63:0] _2237;
  wire [63:0] _2236;
  wire [63:0] _2235;
  wire [63:0] _2234;
  wire [63:0] _2233;
  wire [63:0] _2232;
  wire [31:0] _2231;
  wire [63:0] _2230;
  wire [63:0] _2229;
  wire [63:0] _2228;
  wire [63:0] _2227;
  wire [63:0] _2226;
  wire [31:0] _2225;
  wire [63:0] _2224;
  wire [63:0] _2223;
  wire [63:0] _2222;
  wire [63:0] _2221;
  wire [63:0] _2220;
  wire [63:0] _2219;
  wire [63:0] _2218;
  wire [63:0] _2217;
  wire [63:0] _2216;
  wire [63:0] _2215;
  wire [63:0] _2214;
  wire [31:0] _2213;
  wire [63:0] _2212;
  wire [63:0] _2211;
  wire [63:0] _2210;
  wire [63:0] _2209;
  wire [63:0] _2208;
  wire [31:0] _2207;
  wire [63:0] _2206;
  wire [63:0] _2205;
  wire [63:0] _2204;
  wire [63:0] _2203;
  wire [63:0] _2202;
  wire [63:0] _2201;
  wire [63:0] _2200;
  wire [63:0] _2199;
  wire [63:0] _2198;
  wire [31:0] _2197;
  wire [63:0] _2196;
  wire [63:0] _2195;
  wire [63:0] _2194;
  wire [63:0] _2193;
  wire [63:0] _2192;
  wire [31:0] _2191;
  wire [63:0] _2190;
  wire [63:0] _2189;
  wire [63:0] _2188;
  wire [63:0] _2187;
  wire [31:0] _2186;
  wire [63:0] _2185;
  wire [63:0] _2184;
  wire [63:0] _2183;
  wire [0:0] ifout2288;
  wire [63:0] _2182;
  wire [63:0] _2181;
  wire [63:0] _2180;
  wire [63:0] _2179;
  wire [63:0] _2178;
  wire [63:0] _2177;
  wire [7:0] _2572;
  wire [63:0] _2176;
  wire [63:0] _2175;
  wire [31:0] n_idx_2571;
  wire [31:0] _2174;
  wire [63:0] _2173;
  wire [63:0] _2172;
  wire [63:0] _2171;
  wire [63:0] _2170;
  wire [63:0] _2169;
  wire [63:0] _2168;
  wire [63:0] _2167;
  wire [63:0] _2166;
  wire [63:0] _2165;
  wire [63:0] _2164;
  wire [63:0] _2163;
  wire [63:0] _2162;
  wire [31:0] _2161;
  wire [63:0] _2160;
  wire [63:0] _2159;
  wire [63:0] _2158;
  wire [63:0] _2157;
  wire [63:0] _2156;
  wire [31:0] _2155;
  wire [63:0] _2154;
  wire [63:0] _2153;
  wire [63:0] _2152;
  wire [63:0] _2151;
  wire [63:0] _2150;
  wire [63:0] _2149;
  wire [63:0] _2148;
  wire [63:0] _2147;
  wire [63:0] _2146;
  wire [31:0] _2145;
  wire [63:0] _2144;
  wire [63:0] _2143;
  wire [63:0] _2142;
  wire [63:0] _2141;
  wire [63:0] _2140;
  wire [31:0] _2139;
  wire [63:0] _2138;
  wire [63:0] _2137;
  wire [63:0] _2136;
  wire [63:0] _2135;
  wire [63:0] _2134;
  wire [63:0] _2133;
  wire [63:0] _2132;
  wire [63:0] _2131;
  wire [63:0] _2130;
  wire [63:0] _2129;
  wire [63:0] _2128;
  wire [31:0] _2127;
  wire [63:0] _2126;
  wire [63:0] _2125;
  wire [63:0] _2124;
  wire [63:0] _2123;
  wire [63:0] _2122;
  wire [31:0] _2121;
  wire [63:0] _2120;
  wire [63:0] _2119;
  wire [63:0] _2118;
  wire [63:0] _2117;
  wire [63:0] _2116;
  wire [63:0] _2115;
  wire [63:0] _2114;
  wire [63:0] _2113;
  wire [63:0] _2112;
  wire [31:0] _2111;
  wire [63:0] _2110;
  wire [63:0] _2109;
  wire [63:0] _2108;
  wire [63:0] _2107;
  wire [63:0] _2106;
  wire [31:0] _2105;
  wire [63:0] _2104;
  wire [63:0] _2103;
  wire [63:0] _2102;
  wire [63:0] _2101;
  wire [31:0] _2100;
  wire [63:0] _2099;
  wire [63:0] _2098;
  wire [63:0] _2097;
  wire [0:0] ifout2199;
  wire [63:0] _2096;
  wire [63:0] _2095;
  wire [63:0] _2094;
  wire [63:0] _2093;
  wire [63:0] _2092;
  wire [63:0] _2091;
  wire [7:0] _2582;
  wire [63:0] _2090;
  wire [63:0] _2089;
  wire [31:0] n_idx_2581;
  wire [31:0] _2088;
  wire [63:0] _2087;
  wire [63:0] _2086;
  wire [63:0] _2085;
  wire [63:0] _2084;
  wire [63:0] _2083;
  wire [63:0] _2082;
  wire [63:0] _2081;
  wire [63:0] _2080;
  wire [63:0] _2079;
  wire [63:0] _2078;
  wire [63:0] _2077;
  wire [63:0] _2076;
  wire [31:0] _2075;
  wire [63:0] _2074;
  wire [63:0] _2073;
  wire [63:0] _2072;
  wire [63:0] _2071;
  wire [63:0] _2070;
  wire [31:0] _2069;
  wire [63:0] _2068;
  wire [63:0] _2067;
  wire [63:0] _2066;
  wire [63:0] _2065;
  wire [63:0] _2064;
  wire [63:0] _2063;
  wire [63:0] _2062;
  wire [63:0] _2061;
  wire [63:0] _2060;
  wire [31:0] _2059;
  wire [63:0] _2058;
  wire [63:0] _2057;
  wire [63:0] _2056;
  wire [63:0] _2055;
  wire [63:0] _2054;
  wire [31:0] _2053;
  wire [63:0] _2052;
  wire [63:0] _2051;
  wire [63:0] _2050;
  wire [63:0] _2049;
  wire [63:0] _2048;
  wire [63:0] _2047;
  wire [63:0] _2046;
  wire [63:0] _2045;
  wire [63:0] _2044;
  wire [63:0] _2043;
  wire [63:0] _2042;
  wire [31:0] _2041;
  wire [63:0] _2040;
  wire [63:0] _2039;
  wire [63:0] _2038;
  wire [63:0] _2037;
  wire [63:0] _2036;
  wire [31:0] _2035;
  wire [63:0] _2034;
  wire [63:0] _2033;
  wire [63:0] _2032;
  wire [63:0] _2031;
  wire [63:0] _2030;
  wire [63:0] _2029;
  wire [63:0] _2028;
  wire [63:0] _2027;
  wire [63:0] _2026;
  wire [31:0] _2025;
  wire [63:0] _2024;
  wire [63:0] _2023;
  wire [63:0] _2022;
  wire [63:0] _2021;
  wire [63:0] _2020;
  wire [31:0] _2019;
  wire [63:0] _2018;
  wire [63:0] _2017;
  wire [63:0] _2016;
  wire [63:0] _2015;
  wire [31:0] _2014;
  wire [63:0] _2013;
  wire [63:0] _2012;
  wire [63:0] _2011;
  wire [0:0] ifout2110;
  wire [63:0] _2010;
  wire [63:0] _2009;
  wire [63:0] _2008;
  wire [63:0] _2007;
  wire [63:0] _2006;
  wire [63:0] _2005;
  wire [7:0] _2592;
  wire [63:0] _2004;
  wire [63:0] _2003;
  wire [31:0] n_idx_2591;
  wire [31:0] _2002;
  wire [63:0] _2001;
  wire [63:0] _2000;
  wire [63:0] _1999;
  wire [63:0] _1998;
  wire [63:0] _1997;
  wire [63:0] _1996;
  wire [63:0] _1995;
  wire [63:0] _1994;
  wire [63:0] _1993;
  wire [63:0] _1992;
  wire [63:0] _1991;
  wire [63:0] _1990;
  wire [31:0] _1989;
  wire [63:0] _1988;
  wire [63:0] _1987;
  wire [63:0] _1986;
  wire [63:0] _1985;
  wire [63:0] _1984;
  wire [31:0] _1983;
  wire [63:0] _1982;
  wire [63:0] _1981;
  wire [63:0] _1980;
  wire [63:0] _1979;
  wire [63:0] _1978;
  wire [63:0] _1977;
  wire [63:0] _1976;
  wire [63:0] _1975;
  wire [63:0] _1974;
  wire [31:0] _1973;
  wire [63:0] _1972;
  wire [63:0] _1971;
  wire [63:0] _1970;
  wire [63:0] _1969;
  wire [63:0] _1968;
  wire [31:0] _1967;
  wire [63:0] _1966;
  wire [63:0] _1965;
  wire [63:0] _1964;
  wire [63:0] _1963;
  wire [63:0] _1962;
  wire [63:0] _1961;
  wire [63:0] _1960;
  wire [63:0] _1959;
  wire [63:0] _1958;
  wire [63:0] _1957;
  wire [63:0] _1956;
  wire [31:0] _1955;
  wire [63:0] _1954;
  wire [63:0] _1953;
  wire [63:0] _1952;
  wire [63:0] _1951;
  wire [63:0] _1950;
  wire [31:0] _1949;
  wire [63:0] _1948;
  wire [63:0] _1947;
  wire [63:0] _1946;
  wire [63:0] _1945;
  wire [63:0] _1944;
  wire [63:0] _1943;
  wire [63:0] _1942;
  wire [63:0] _1941;
  wire [63:0] _1940;
  wire [31:0] _1939;
  wire [63:0] _1938;
  wire [63:0] _1937;
  wire [63:0] _1936;
  wire [63:0] _1935;
  wire [63:0] _1934;
  wire [31:0] _1933;
  wire [63:0] _1932;
  wire [63:0] _1931;
  wire [63:0] _1930;
  wire [63:0] _1929;
  wire [31:0] _1928;
  wire [63:0] _1927;
  wire [63:0] _1926;
  wire [63:0] _1925;
  wire [0:0] ifout2021;
  wire [63:0] _1924;
  wire [63:0] _1923;
  wire [63:0] _1922;
  wire [63:0] _1921;
  wire [63:0] _1920;
  wire [63:0] _1919;
  wire [7:0] _2603;
  wire [63:0] _1918;
  wire [63:0] _1917;
  wire [31:0] n_idx_2602;
  wire [31:0] _1916;
  wire [63:0] _1915;
  wire [63:0] _1914;
  wire [63:0] _1913;
  wire [63:0] _1912;
  wire [63:0] _1911;
  wire [63:0] _1910;
  wire [63:0] _1909;
  wire [63:0] _1908;
  wire [63:0] _1907;
  wire [63:0] _1906;
  wire [63:0] _1905;
  wire [63:0] _1904;
  wire [31:0] _1903;
  wire [63:0] _1902;
  wire [63:0] _1901;
  wire [63:0] _1900;
  wire [63:0] _1899;
  wire [63:0] _1898;
  wire [31:0] _1897;
  wire [63:0] _1896;
  wire [63:0] _1895;
  wire [63:0] _1894;
  wire [63:0] _1893;
  wire [63:0] _1892;
  wire [63:0] _1891;
  wire [63:0] _1890;
  wire [63:0] _1889;
  wire [63:0] _1888;
  wire [31:0] _1887;
  wire [63:0] _1886;
  wire [63:0] _1885;
  wire [63:0] _1884;
  wire [63:0] _1883;
  wire [63:0] _1882;
  wire [31:0] _1881;
  wire [63:0] _1880;
  wire [63:0] _1879;
  wire [63:0] _1878;
  wire [63:0] _1877;
  wire [63:0] _1876;
  wire [63:0] _1875;
  wire [63:0] _1874;
  wire [63:0] _1873;
  wire [63:0] _1872;
  wire [63:0] _1871;
  wire [63:0] _1870;
  wire [31:0] _1869;
  wire [63:0] _1868;
  wire [63:0] _1867;
  wire [63:0] _1866;
  wire [63:0] _1865;
  wire [63:0] _1864;
  wire [31:0] _1863;
  wire [63:0] _1862;
  wire [63:0] _1861;
  wire [63:0] _1860;
  wire [63:0] _1859;
  wire [63:0] _1858;
  wire [63:0] _1857;
  wire [63:0] _1856;
  wire [63:0] _1855;
  wire [63:0] _1854;
  wire [31:0] _1853;
  wire [63:0] _1852;
  wire [63:0] _1851;
  wire [63:0] _1850;
  wire [63:0] _1849;
  wire [63:0] _1848;
  wire [31:0] _1847;
  wire [63:0] _1846;
  wire [63:0] _1845;
  wire [63:0] _1844;
  wire [63:0] _1843;
  wire [31:0] _1842;
  wire [63:0] _1841;
  wire [63:0] _1840;
  wire [63:0] _1839;
  wire [0:0] ifout1932;
  wire [63:0] _1838;
  wire [63:0] _1837;
  wire [63:0] _1836;
  wire [63:0] _1835;
  wire [63:0] _1834;
  wire [63:0] _1833;
  wire [7:0] _2613;
  wire [63:0] _1832;
  wire [63:0] _1831;
  wire [31:0] n_idx_2612;
  wire [31:0] _1830;
  wire [63:0] _1829;
  wire [63:0] _1828;
  wire [63:0] _1827;
  wire [63:0] _1826;
  wire [63:0] _1825;
  wire [63:0] _1824;
  wire [63:0] _1823;
  wire [63:0] _1822;
  wire [63:0] _1821;
  wire [63:0] _1820;
  wire [63:0] _1819;
  wire [63:0] _1818;
  wire [31:0] _1817;
  wire [63:0] _1816;
  wire [63:0] _1815;
  wire [63:0] _1814;
  wire [63:0] _1813;
  wire [63:0] _1812;
  wire [31:0] _1811;
  wire [63:0] _1810;
  wire [63:0] _1809;
  wire [63:0] _1808;
  wire [63:0] _1807;
  wire [63:0] _1806;
  wire [63:0] _1805;
  wire [63:0] _1804;
  wire [63:0] _1803;
  wire [63:0] _1802;
  wire [31:0] _1801;
  wire [63:0] _1800;
  wire [63:0] _1799;
  wire [63:0] _1798;
  wire [63:0] _1797;
  wire [63:0] _1796;
  wire [31:0] _1795;
  wire [63:0] _1794;
  wire [63:0] _1793;
  wire [63:0] _1792;
  wire [63:0] _1791;
  wire [63:0] _1790;
  wire [63:0] _1789;
  wire [63:0] _1788;
  wire [63:0] _1787;
  wire [63:0] _1786;
  wire [63:0] _1785;
  wire [63:0] _1784;
  wire [31:0] _1783;
  wire [63:0] _1782;
  wire [63:0] _1781;
  wire [63:0] _1780;
  wire [63:0] _1779;
  wire [63:0] _1778;
  wire [31:0] _1777;
  wire [63:0] _1776;
  wire [63:0] _1775;
  wire [63:0] _1774;
  wire [63:0] _1773;
  wire [63:0] _1772;
  wire [63:0] _1771;
  wire [63:0] _1770;
  wire [63:0] _1769;
  wire [63:0] _1768;
  wire [31:0] _1767;
  wire [63:0] _1766;
  wire [63:0] _1765;
  wire [63:0] _1764;
  wire [63:0] _1763;
  wire [63:0] _1762;
  wire [31:0] _1761;
  wire [63:0] _1760;
  wire [63:0] _1759;
  wire [63:0] _1758;
  wire [63:0] _1757;
  wire [31:0] _1756;
  wire [63:0] _1755;
  wire [63:0] _1754;
  wire [63:0] _1753;
  wire [0:0] ifout1843;
  wire [63:0] _1752;
  wire [63:0] _1751;
  wire [63:0] _1750;
  wire [63:0] _1749;
  wire [63:0] _1748;
  wire [63:0] _1747;
  wire [7:0] _2623;
  wire [63:0] _1746;
  wire [63:0] _1745;
  wire [31:0] n_idx_2622;
  wire [31:0] _1744;
  wire [63:0] _1743;
  wire [63:0] _1742;
  wire [63:0] _1741;
  wire [63:0] _1740;
  wire [63:0] _1739;
  wire [63:0] _1738;
  wire [63:0] _1737;
  wire [63:0] _1736;
  wire [63:0] _1735;
  wire [63:0] _1734;
  wire [63:0] _1733;
  wire [63:0] _1732;
  wire [31:0] _1731;
  wire [63:0] _1730;
  wire [63:0] _1729;
  wire [63:0] _1728;
  wire [63:0] _1727;
  wire [63:0] _1726;
  wire [31:0] _1725;
  wire [63:0] _1724;
  wire [63:0] _1723;
  wire [63:0] _1722;
  wire [63:0] _1721;
  wire [63:0] _1720;
  wire [63:0] _1719;
  wire [63:0] _1718;
  wire [63:0] _1717;
  wire [63:0] _1716;
  wire [31:0] _1715;
  wire [63:0] _1714;
  wire [63:0] _1713;
  wire [63:0] _1712;
  wire [63:0] _1711;
  wire [63:0] _1710;
  wire [31:0] _1709;
  wire [63:0] _1708;
  wire [63:0] _1707;
  wire [63:0] _1706;
  wire [63:0] _1705;
  wire [63:0] _1704;
  wire [63:0] _1703;
  wire [63:0] _1702;
  wire [63:0] _1701;
  wire [63:0] _1700;
  wire [63:0] _1699;
  wire [63:0] _1698;
  wire [31:0] _1697;
  wire [63:0] _1696;
  wire [63:0] _1695;
  wire [63:0] _1694;
  wire [63:0] _1693;
  wire [63:0] _1692;
  wire [31:0] _1691;
  wire [63:0] _1690;
  wire [63:0] _1689;
  wire [63:0] _1688;
  wire [63:0] _1687;
  wire [63:0] _1686;
  wire [63:0] _1685;
  wire [63:0] _1684;
  wire [63:0] _1683;
  wire [63:0] _1682;
  wire [31:0] _1681;
  wire [63:0] _1680;
  wire [63:0] _1679;
  wire [63:0] _1678;
  wire [63:0] _1677;
  wire [63:0] _1676;
  wire [31:0] _1675;
  wire [63:0] _1674;
  wire [63:0] _1673;
  wire [63:0] _1672;
  wire [63:0] _1671;
  wire [31:0] _1670;
  wire [63:0] _1669;
  wire [63:0] _1668;
  wire [63:0] _1667;
  wire [0:0] ifout1754;
  wire [63:0] _1666;
  wire [63:0] _1665;
  wire [63:0] _1664;
  wire [63:0] _1663;
  wire [63:0] _1662;
  wire [63:0] _1661;
  wire [7:0] _2633;
  wire [63:0] _1660;
  wire [63:0] _1659;
  wire [31:0] n_idx_2632;
  wire [31:0] _1658;
  wire [63:0] _1657;
  wire [63:0] _1656;
  wire [63:0] _1655;
  wire [63:0] _1654;
  wire [63:0] _1653;
  wire [63:0] _1652;
  wire [63:0] _1651;
  wire [63:0] _1650;
  wire [63:0] _1649;
  wire [63:0] _1648;
  wire [63:0] _1647;
  wire [63:0] _1646;
  wire [31:0] _1645;
  wire [63:0] _1644;
  wire [63:0] _1643;
  wire [63:0] _1642;
  wire [63:0] _1641;
  wire [63:0] _1640;
  wire [31:0] _1639;
  wire [63:0] _1638;
  wire [63:0] _1637;
  wire [63:0] _1636;
  wire [63:0] _1635;
  wire [63:0] _1634;
  wire [63:0] _1633;
  wire [63:0] _1632;
  wire [63:0] _1631;
  wire [63:0] _1630;
  wire [31:0] _1629;
  wire [63:0] _1628;
  wire [63:0] _1627;
  wire [63:0] _1626;
  wire [63:0] _1625;
  wire [63:0] _1624;
  wire [31:0] _1623;
  wire [63:0] _1622;
  wire [63:0] _1621;
  wire [63:0] _1620;
  wire [63:0] _1619;
  wire [63:0] _1618;
  wire [63:0] _1617;
  wire [63:0] _1616;
  wire [63:0] _1615;
  wire [63:0] _1614;
  wire [63:0] _1613;
  wire [63:0] _1612;
  wire [31:0] _1611;
  wire [63:0] _1610;
  wire [63:0] _1609;
  wire [63:0] _1608;
  wire [63:0] _1607;
  wire [63:0] _1606;
  wire [31:0] _1605;
  wire [63:0] _1604;
  wire [63:0] _1603;
  wire [63:0] _1602;
  wire [63:0] _1601;
  wire [63:0] _1600;
  wire [63:0] _1599;
  wire [63:0] _1598;
  wire [63:0] _1597;
  wire [63:0] _1596;
  wire [31:0] _1595;
  wire [63:0] _1594;
  wire [63:0] _1593;
  wire [63:0] _1592;
  wire [63:0] _1591;
  wire [63:0] _1590;
  wire [31:0] _1589;
  wire [63:0] _1588;
  wire [63:0] _1587;
  wire [63:0] _1586;
  wire [63:0] _1585;
  wire [31:0] _1584;
  wire [63:0] _1583;
  wire [63:0] _1582;
  wire [63:0] _1581;
  wire [0:0] ifout1665;
  wire [63:0] _1580;
  wire [63:0] _1579;
  wire [63:0] _1578;
  wire [63:0] _1577;
  wire [63:0] _1576;
  wire [63:0] _1575;
  wire [7:0] _2643;
  wire [63:0] _1574;
  wire [63:0] _1573;
  wire [31:0] n_idx_2642;
  wire [31:0] _1572;
  wire [63:0] _1571;
  wire [63:0] _1570;
  wire [63:0] _1569;
  wire [63:0] _1568;
  wire [63:0] _1567;
  wire [63:0] _1566;
  wire [63:0] _1565;
  wire [63:0] _1564;
  wire [63:0] _1563;
  wire [63:0] _1562;
  wire [63:0] _1561;
  wire [63:0] _1560;
  wire [31:0] _1559;
  wire [63:0] _1558;
  wire [63:0] _1557;
  wire [63:0] _1556;
  wire [63:0] _1555;
  wire [63:0] _1554;
  wire [31:0] _1553;
  wire [63:0] _1552;
  wire [63:0] _1551;
  wire [63:0] _1550;
  wire [63:0] _1549;
  wire [63:0] _1548;
  wire [63:0] _1547;
  wire [63:0] _1546;
  wire [63:0] _1545;
  wire [63:0] _1544;
  wire [31:0] _1543;
  wire [63:0] _1542;
  wire [63:0] _1541;
  wire [63:0] _1540;
  wire [63:0] _1539;
  wire [63:0] _1538;
  wire [31:0] _1537;
  wire [63:0] _1536;
  wire [63:0] _1535;
  wire [63:0] _1534;
  wire [63:0] _1533;
  wire [63:0] _1532;
  wire [63:0] _1531;
  wire [63:0] _1530;
  wire [63:0] _1529;
  wire [63:0] _1528;
  wire [63:0] _1527;
  wire [63:0] _1526;
  wire [31:0] _1525;
  wire [63:0] _1524;
  wire [63:0] _1523;
  wire [63:0] _1522;
  wire [63:0] _1521;
  wire [63:0] _1520;
  wire [31:0] _1519;
  wire [63:0] _1518;
  wire [63:0] _1517;
  wire [63:0] _1516;
  wire [63:0] _1515;
  wire [63:0] _1514;
  wire [63:0] _1513;
  wire [63:0] _1512;
  wire [63:0] _1511;
  wire [63:0] _1510;
  wire [31:0] _1509;
  wire [63:0] _1508;
  wire [63:0] _1507;
  wire [63:0] _1506;
  wire [63:0] _1505;
  wire [63:0] _1504;
  wire [31:0] _1503;
  wire [63:0] _1502;
  wire [63:0] _1501;
  wire [63:0] _1500;
  wire [63:0] _1499;
  wire [31:0] _1498;
  wire [63:0] _1497;
  wire [63:0] _1496;
  wire [63:0] _1495;
  wire [0:0] ifout1576;
  wire [63:0] _1494;
  wire [63:0] _1493;
  wire [63:0] _1492;
  wire [63:0] _1491;
  wire [63:0] _1490;
  wire [63:0] _1489;
  wire [7:0] _2653;
  wire [63:0] _1488;
  wire [63:0] _1487;
  wire [31:0] n_idx_2652;
  wire [31:0] _1486;
  wire [63:0] _1485;
  wire [63:0] _1484;
  wire [63:0] _1483;
  wire [63:0] _1482;
  wire [63:0] _1481;
  wire [63:0] _1480;
  wire [63:0] _1479;
  wire [63:0] _1478;
  wire [63:0] _1477;
  wire [63:0] _1476;
  wire [63:0] _1475;
  wire [63:0] _1474;
  wire [31:0] _1473;
  wire [63:0] _1472;
  wire [63:0] _1471;
  wire [63:0] _1470;
  wire [63:0] _1469;
  wire [63:0] _1468;
  wire [31:0] _1467;
  wire [63:0] _1466;
  wire [63:0] _1465;
  wire [63:0] _1464;
  wire [63:0] _1463;
  wire [63:0] _1462;
  wire [63:0] _1461;
  wire [63:0] _1460;
  wire [63:0] _1459;
  wire [63:0] _1458;
  wire [31:0] _1457;
  wire [63:0] _1456;
  wire [63:0] _1455;
  wire [63:0] _1454;
  wire [63:0] _1453;
  wire [63:0] _1452;
  wire [31:0] _1451;
  wire [63:0] _1450;
  wire [63:0] _1449;
  wire [63:0] _1448;
  wire [63:0] _1447;
  wire [63:0] _1446;
  wire [63:0] _1445;
  wire [63:0] _1444;
  wire [63:0] _1443;
  wire [63:0] _1442;
  wire [63:0] _1441;
  wire [63:0] _1440;
  wire [31:0] _1439;
  wire [63:0] _1438;
  wire [63:0] _1437;
  wire [63:0] _1436;
  wire [63:0] _1435;
  wire [63:0] _1434;
  wire [31:0] _1433;
  wire [63:0] _1432;
  wire [63:0] _1431;
  wire [63:0] _1430;
  wire [63:0] _1429;
  wire [63:0] _1428;
  wire [63:0] _1427;
  wire [63:0] _1426;
  wire [63:0] _1425;
  wire [63:0] _1424;
  wire [31:0] _1423;
  wire [63:0] _1422;
  wire [63:0] _1421;
  wire [63:0] _1420;
  wire [63:0] _1419;
  wire [63:0] _1418;
  wire [31:0] _1417;
  wire [63:0] _1416;
  wire [63:0] _1415;
  wire [63:0] _1414;
  wire [63:0] _1413;
  wire [31:0] _1412;
  wire [63:0] _1411;
  wire [63:0] _1410;
  wire [63:0] _1409;
  wire [0:0] ifout1487;
  wire [63:0] _1408;
  wire [63:0] _1407;
  wire [63:0] _1406;
  wire [63:0] _1405;
  wire [63:0] _1404;
  wire [63:0] _1403;
  wire [7:0] _2663;
  wire [63:0] _1402;
  wire [63:0] _1401;
  wire [31:0] n_idx_2662;
  wire [31:0] _1400;
  wire [63:0] _1399;
  wire [63:0] _1398;
  wire [63:0] _1397;
  wire [63:0] _1396;
  wire [63:0] _1395;
  wire [63:0] _1394;
  wire [63:0] _1393;
  wire [63:0] _1392;
  wire [63:0] _1391;
  wire [63:0] _1390;
  wire [63:0] _1389;
  wire [63:0] _1388;
  wire [31:0] _1387;
  wire [63:0] _1386;
  wire [63:0] _1385;
  wire [63:0] _1384;
  wire [63:0] _1383;
  wire [63:0] _1382;
  wire [31:0] _1381;
  wire [63:0] _1380;
  wire [63:0] _1379;
  wire [63:0] _1378;
  wire [63:0] _1377;
  wire [63:0] _1376;
  wire [63:0] _1375;
  wire [63:0] _1374;
  wire [63:0] _1373;
  wire [63:0] _1372;
  wire [31:0] _1371;
  wire [63:0] _1370;
  wire [63:0] _1369;
  wire [63:0] _1368;
  wire [63:0] _1367;
  wire [63:0] _1366;
  wire [31:0] _1365;
  wire [63:0] _1364;
  wire [63:0] _1363;
  wire [63:0] _1362;
  wire [63:0] _1361;
  wire [63:0] _1360;
  wire [63:0] _1359;
  wire [63:0] _1358;
  wire [63:0] _1357;
  wire [63:0] _1356;
  wire [63:0] _1355;
  wire [63:0] _1354;
  wire [31:0] _1353;
  wire [63:0] _1352;
  wire [63:0] _1351;
  wire [63:0] _1350;
  wire [63:0] _1349;
  wire [63:0] _1348;
  wire [31:0] _1347;
  wire [63:0] _1346;
  wire [63:0] _1345;
  wire [63:0] _1344;
  wire [63:0] _1343;
  wire [63:0] _1342;
  wire [63:0] _1341;
  wire [63:0] _1340;
  wire [63:0] _1339;
  wire [63:0] _1338;
  wire [31:0] _1337;
  wire [63:0] _1336;
  wire [63:0] _1335;
  wire [63:0] _1334;
  wire [63:0] _1333;
  wire [63:0] _1332;
  wire [31:0] _1331;
  wire [63:0] _1330;
  wire [63:0] _1329;
  wire [63:0] _1328;
  wire [63:0] _1327;
  wire [31:0] _1326;
  wire [63:0] _1325;
  wire [63:0] _1324;
  wire [63:0] _1323;
  wire [0:0] ifout1398;
  wire [63:0] _1322;
  wire [63:0] _1321;
  wire [63:0] _1320;
  wire [63:0] _1319;
  wire [63:0] _1318;
  wire [63:0] _1317;
  wire [7:0] _2672;
  wire [63:0] _1316;
  wire [63:0] _1315;
  wire [31:0] n_idx_2671;
  wire [31:0] _1314;
  wire [63:0] _1313;
  wire [63:0] _1312;
  wire [63:0] _1311;
  wire [63:0] _1310;
  wire [63:0] _1309;
  wire [63:0] _1308;
  wire [63:0] _1307;
  wire [63:0] _1306;
  wire [63:0] _1305;
  wire [63:0] _1304;
  wire [63:0] _1303;
  wire [63:0] _1302;
  wire [31:0] _1301;
  wire [63:0] _1300;
  wire [63:0] _1299;
  wire [63:0] _1298;
  wire [63:0] _1297;
  wire [63:0] _1296;
  wire [31:0] _1295;
  wire [63:0] _1294;
  wire [63:0] _1293;
  wire [63:0] _1292;
  wire [63:0] _1291;
  wire [63:0] _1290;
  wire [63:0] _1289;
  wire [63:0] _1288;
  wire [63:0] _1287;
  wire [63:0] _1286;
  wire [31:0] _1285;
  wire [63:0] _1284;
  wire [63:0] _1283;
  wire [63:0] _1282;
  wire [63:0] _1281;
  wire [63:0] _1280;
  wire [31:0] _1279;
  wire [63:0] _1278;
  wire [63:0] _1277;
  wire [63:0] _1276;
  wire [63:0] _1275;
  wire [63:0] _1274;
  wire [63:0] _1273;
  wire [63:0] _1272;
  wire [63:0] _1271;
  wire [63:0] _1270;
  wire [63:0] _1269;
  wire [63:0] _1268;
  wire [31:0] _1267;
  wire [63:0] _1266;
  wire [63:0] _1265;
  wire [63:0] _1264;
  wire [63:0] _1263;
  wire [63:0] _1262;
  wire [31:0] _1261;
  wire [63:0] _1260;
  wire [63:0] _1259;
  wire [63:0] _1258;
  wire [63:0] _1257;
  wire [63:0] _1256;
  wire [63:0] _1255;
  wire [63:0] _1254;
  wire [63:0] _1253;
  wire [63:0] _1252;
  wire [31:0] _1251;
  wire [63:0] _1250;
  wire [63:0] _1249;
  wire [63:0] _1248;
  wire [63:0] _1247;
  wire [63:0] _1246;
  wire [31:0] _1245;
  wire [63:0] _1244;
  wire [63:0] _1243;
  wire [63:0] _1242;
  wire [63:0] _1241;
  wire [31:0] _1240;
  wire [63:0] _1239;
  wire [63:0] _1238;
  wire [63:0] _1237;
  wire [0:0] ifout1309;
  wire [63:0] _1236;
  wire [63:0] _1235;
  wire [63:0] _1234;
  wire [63:0] _1233;
  wire [63:0] _1232;
  wire [63:0] _1231;
  wire [31:0] off_2668;
  wire [31:0] idx_2667;
  wire [31:0] idx_sail_2666;
  wire [31:0] _1230;
  wire [31:0] _1229;
  wire [31:0] _1228;
  wire [31:0] ck_idx_2665;
  wire [31:0] _1227;
  wire [63:0] _1226;
  wire [63:0] _1225;
  wire [63:0] _1224;
  wire [63:0] _1223;
  wire [63:0] _1222;
  wire [63:0] _1221;
  wire [63:0] _1220;
  wire [63:0] _1219;
  wire [63:0] _1218;
  wire [63:0] _1217;
  wire [63:0] _1216;
  wire [63:0] _1215;
  wire [31:0] _1214;
  wire [63:0] _1213;
  wire [63:0] _1212;
  wire [63:0] _1211;
  wire [63:0] _1210;
  wire [63:0] _1209;
  wire [31:0] _1208;
  wire [63:0] _1207;
  wire [63:0] _1206;
  wire [63:0] _1205;
  wire [63:0] _1204;
  wire [63:0] _1203;
  wire [63:0] _1202;
  wire [63:0] _1201;
  wire [63:0] _1200;
  wire [63:0] _1199;
  wire [31:0] _1198;
  wire [63:0] _1197;
  wire [63:0] _1196;
  wire [63:0] _1195;
  wire [63:0] _1194;
  wire [63:0] _1193;
  wire [31:0] _1192;
  wire [63:0] _1191;
  wire [63:0] _1190;
  wire [63:0] _1189;
  wire [63:0] _1188;
  wire [63:0] _1187;
  wire [63:0] _1186;
  wire [63:0] _1185;
  wire [63:0] _1184;
  wire [63:0] _1183;
  wire [63:0] _1182;
  wire [63:0] _1181;
  wire [31:0] _1180;
  wire [63:0] _1179;
  wire [63:0] _1178;
  wire [63:0] _1177;
  wire [63:0] _1176;
  wire [63:0] _1175;
  wire [31:0] _1174;
  wire [63:0] _1173;
  wire [63:0] _1172;
  wire [63:0] _1171;
  wire [63:0] _1170;
  wire [63:0] _1169;
  wire [63:0] _1168;
  wire [63:0] _1167;
  wire [63:0] _1166;
  wire [63:0] _1165;
  wire [31:0] _1164;
  wire [63:0] _1163;
  wire [63:0] _1162;
  wire [63:0] _1161;
  wire [63:0] _1160;
  wire [63:0] _1159;
  wire [31:0] _1158;
  wire [63:0] _1157;
  wire [63:0] _1156;
  wire [63:0] _1155;
  wire [63:0] _1154;
  wire [31:0] _1153;
  wire [63:0] _1152;
  wire [63:0] _1151;
  wire [63:0] _1150;
  wire [0:0] ifout1217;
  wire [63:0] _1149;
  wire [63:0] _1148;
  wire [63:0] _1147;
  wire [63:0] _1146;
  wire [63:0] _1145;
  wire [63:0] _1144;
  wire [31:0] off_2658;
  wire [31:0] idx_2657;
  wire [31:0] idx_sail_2656;
  wire [31:0] _1143;
  wire [31:0] _1142;
  wire [63:0] _1141;
  wire [31:0] _1140;
  wire [31:0] ck_idx_2655;
  wire [31:0] _1139;
  wire [63:0] _1138;
  wire [63:0] _1137;
  wire [63:0] _1136;
  wire [63:0] _1135;
  wire [63:0] _1134;
  wire [63:0] _1133;
  wire [63:0] _1132;
  wire [63:0] _1131;
  wire [63:0] _1130;
  wire [63:0] _1129;
  wire [63:0] _1128;
  wire [63:0] _1127;
  wire [31:0] _1126;
  wire [63:0] _1125;
  wire [63:0] _1124;
  wire [63:0] _1123;
  wire [63:0] _1122;
  wire [63:0] _1121;
  wire [31:0] _1120;
  wire [63:0] _1119;
  wire [63:0] _1118;
  wire [63:0] _1117;
  wire [63:0] _1116;
  wire [63:0] _1115;
  wire [63:0] _1114;
  wire [63:0] _1113;
  wire [63:0] _1112;
  wire [63:0] _1111;
  wire [31:0] _1110;
  wire [63:0] _1109;
  wire [63:0] _1108;
  wire [63:0] _1107;
  wire [63:0] _1106;
  wire [63:0] _1105;
  wire [31:0] _1104;
  wire [63:0] _1103;
  wire [63:0] _1102;
  wire [63:0] _1101;
  wire [63:0] _1100;
  wire [63:0] _1099;
  wire [63:0] _1098;
  wire [63:0] _1097;
  wire [63:0] _1096;
  wire [63:0] _1095;
  wire [63:0] _1094;
  wire [63:0] _1093;
  wire [31:0] _1092;
  wire [63:0] _1091;
  wire [63:0] _1090;
  wire [63:0] _1089;
  wire [63:0] _1088;
  wire [63:0] _1087;
  wire [31:0] _1086;
  wire [63:0] _1085;
  wire [63:0] _1084;
  wire [63:0] _1083;
  wire [63:0] _1082;
  wire [63:0] _1081;
  wire [63:0] _1080;
  wire [63:0] _1079;
  wire [63:0] _1078;
  wire [63:0] _1077;
  wire [31:0] _1076;
  wire [63:0] _1075;
  wire [63:0] _1074;
  wire [63:0] _1073;
  wire [63:0] _1072;
  wire [63:0] _1071;
  wire [31:0] _1070;
  wire [63:0] _1069;
  wire [63:0] _1068;
  wire [63:0] _1067;
  wire [63:0] _1066;
  wire [31:0] _1065;
  wire [63:0] _1064;
  wire [63:0] _1063;
  wire [63:0] _1062;
  wire [0:0] ifout1124;
  wire [63:0] _1061;
  wire [63:0] _1060;
  wire [63:0] _1059;
  wire [63:0] _1058;
  wire [63:0] _1057;
  wire [63:0] _1056;
  wire [31:0] off_2648;
  wire [31:0] idx_2647;
  wire [31:0] idx_sail_2646;
  wire [31:0] _1055;
  wire [31:0] _1054;
  wire [63:0] _1053;
  wire [31:0] _1052;
  wire [31:0] ck_idx_2645;
  wire [31:0] _1051;
  wire [63:0] _1050;
  wire [63:0] _1049;
  wire [63:0] _1048;
  wire [63:0] _1047;
  wire [63:0] _1046;
  wire [63:0] _1045;
  wire [63:0] _1044;
  wire [63:0] _1043;
  wire [63:0] _1042;
  wire [63:0] _1041;
  wire [63:0] _1040;
  wire [63:0] _1039;
  wire [31:0] _1038;
  wire [63:0] _1037;
  wire [63:0] _1036;
  wire [63:0] _1035;
  wire [63:0] _1034;
  wire [63:0] _1033;
  wire [31:0] _1032;
  wire [63:0] _1031;
  wire [63:0] _1030;
  wire [63:0] _1029;
  wire [63:0] _1028;
  wire [63:0] _1027;
  wire [63:0] _1026;
  wire [63:0] _1025;
  wire [63:0] _1024;
  wire [63:0] _1023;
  wire [31:0] _1022;
  wire [63:0] _1021;
  wire [63:0] _1020;
  wire [63:0] _1019;
  wire [63:0] _1018;
  wire [63:0] _1017;
  wire [31:0] _1016;
  wire [63:0] _1015;
  wire [63:0] _1014;
  wire [63:0] _1013;
  wire [63:0] _1012;
  wire [63:0] _1011;
  wire [63:0] _1010;
  wire [63:0] _1009;
  wire [63:0] _1008;
  wire [63:0] _1007;
  wire [63:0] _1006;
  wire [63:0] _1005;
  wire [31:0] _1004;
  wire [63:0] _1003;
  wire [63:0] _1002;
  wire [63:0] _1001;
  wire [63:0] _1000;
  wire [63:0] _999;
  wire [31:0] _998;
  wire [63:0] _997;
  wire [63:0] _996;
  wire [63:0] _995;
  wire [63:0] _994;
  wire [63:0] _993;
  wire [63:0] _992;
  wire [63:0] _991;
  wire [63:0] _990;
  wire [63:0] _989;
  wire [31:0] _988;
  wire [63:0] _987;
  wire [63:0] _986;
  wire [63:0] _985;
  wire [63:0] _984;
  wire [63:0] _983;
  wire [31:0] _982;
  wire [63:0] _981;
  wire [63:0] _980;
  wire [63:0] _979;
  wire [63:0] _978;
  wire [31:0] _977;
  wire [63:0] _976;
  wire [63:0] _975;
  wire [63:0] _974;
  wire [0:0] ifout1031;
  wire [63:0] _973;
  wire [63:0] _972;
  wire [63:0] _971;
  wire [63:0] _970;
  wire [63:0] _969;
  wire [63:0] _968;
  wire [31:0] off_2638;
  wire [31:0] idx_2637;
  wire [31:0] idx_sail_2636;
  wire [31:0] _967;
  wire [31:0] _966;
  wire [63:0] _965;
  wire [31:0] _964;
  wire [31:0] ck_idx_2635;
  wire [31:0] _963;
  wire [63:0] _962;
  wire [63:0] _961;
  wire [63:0] _960;
  wire [63:0] _959;
  wire [63:0] _958;
  wire [63:0] _957;
  wire [63:0] _956;
  wire [63:0] _955;
  wire [63:0] _954;
  wire [63:0] _953;
  wire [63:0] _952;
  wire [63:0] _951;
  wire [31:0] _950;
  wire [63:0] _949;
  wire [63:0] _948;
  wire [63:0] _947;
  wire [63:0] _946;
  wire [63:0] _945;
  wire [31:0] _944;
  wire [63:0] _943;
  wire [63:0] _942;
  wire [63:0] _941;
  wire [63:0] _940;
  wire [63:0] _939;
  wire [63:0] _938;
  wire [63:0] _937;
  wire [63:0] _936;
  wire [63:0] _935;
  wire [31:0] _934;
  wire [63:0] _933;
  wire [63:0] _932;
  wire [63:0] _931;
  wire [63:0] _930;
  wire [63:0] _929;
  wire [31:0] _928;
  wire [63:0] _927;
  wire [63:0] _926;
  wire [63:0] _925;
  wire [63:0] _924;
  wire [63:0] _923;
  wire [63:0] _922;
  wire [63:0] _921;
  wire [63:0] _920;
  wire [63:0] _919;
  wire [63:0] _918;
  wire [63:0] _917;
  wire [31:0] _916;
  wire [63:0] _915;
  wire [63:0] _914;
  wire [63:0] _913;
  wire [63:0] _912;
  wire [63:0] _911;
  wire [31:0] _910;
  wire [63:0] _909;
  wire [63:0] _908;
  wire [63:0] _907;
  wire [63:0] _906;
  wire [63:0] _905;
  wire [63:0] _904;
  wire [63:0] _903;
  wire [63:0] _902;
  wire [63:0] _901;
  wire [31:0] _900;
  wire [63:0] _899;
  wire [63:0] _898;
  wire [63:0] _897;
  wire [63:0] _896;
  wire [63:0] _895;
  wire [31:0] _894;
  wire [63:0] _893;
  wire [63:0] _892;
  wire [63:0] _891;
  wire [63:0] _890;
  wire [31:0] _889;
  wire [63:0] _888;
  wire [63:0] _887;
  wire [63:0] _886;
  wire [0:0] ifout938;
  wire [63:0] _885;
  wire [63:0] _884;
  wire [63:0] _883;
  wire [63:0] _882;
  wire [63:0] _881;
  wire [63:0] _880;
  wire [31:0] off_2628;
  wire [31:0] idx_2627;
  wire [31:0] idx_sail_2626;
  wire [31:0] _879;
  wire [31:0] _878;
  wire [63:0] _877;
  wire [31:0] _876;
  wire [31:0] ck_idx_2625;
  wire [31:0] _875;
  wire [63:0] _874;
  wire [63:0] _873;
  wire [63:0] _872;
  wire [63:0] _871;
  wire [63:0] _870;
  wire [63:0] _869;
  wire [63:0] _868;
  wire [63:0] _867;
  wire [63:0] _866;
  wire [63:0] _865;
  wire [63:0] _864;
  wire [63:0] _863;
  wire [31:0] _862;
  wire [63:0] _861;
  wire [63:0] _860;
  wire [63:0] _859;
  wire [63:0] _858;
  wire [63:0] _857;
  wire [31:0] _856;
  wire [63:0] _855;
  wire [63:0] _854;
  wire [63:0] _853;
  wire [63:0] _852;
  wire [63:0] _851;
  wire [63:0] _850;
  wire [63:0] _849;
  wire [63:0] _848;
  wire [63:0] _847;
  wire [31:0] _846;
  wire [63:0] _845;
  wire [63:0] _844;
  wire [63:0] _843;
  wire [63:0] _842;
  wire [63:0] _841;
  wire [31:0] _840;
  wire [63:0] _839;
  wire [63:0] _838;
  wire [63:0] _837;
  wire [63:0] _836;
  wire [63:0] _835;
  wire [63:0] _834;
  wire [63:0] _833;
  wire [63:0] _832;
  wire [63:0] _831;
  wire [63:0] _830;
  wire [63:0] _829;
  wire [31:0] _828;
  wire [63:0] _827;
  wire [63:0] _826;
  wire [63:0] _825;
  wire [63:0] _824;
  wire [63:0] _823;
  wire [31:0] _822;
  wire [63:0] _821;
  wire [63:0] _820;
  wire [63:0] _819;
  wire [63:0] _818;
  wire [63:0] _817;
  wire [63:0] _816;
  wire [63:0] _815;
  wire [63:0] _814;
  wire [63:0] _813;
  wire [31:0] _812;
  wire [63:0] _811;
  wire [63:0] _810;
  wire [63:0] _809;
  wire [63:0] _808;
  wire [63:0] _807;
  wire [31:0] _806;
  wire [63:0] _805;
  wire [63:0] _804;
  wire [63:0] _803;
  wire [63:0] _802;
  wire [31:0] _801;
  wire [63:0] _800;
  wire [63:0] _799;
  wire [63:0] _798;
  wire [0:0] ifout845;
  wire [63:0] _797;
  wire [63:0] _796;
  wire [63:0] _795;
  wire [63:0] _794;
  wire [63:0] _793;
  wire [63:0] _792;
  wire [31:0] off_2618;
  wire [31:0] idx_2617;
  wire [31:0] idx_sail_2616;
  wire [31:0] _791;
  wire [31:0] _790;
  wire [63:0] _789;
  wire [31:0] _788;
  wire [31:0] ck_idx_2615;
  wire [31:0] _787;
  wire [63:0] _786;
  wire [63:0] _785;
  wire [63:0] _784;
  wire [63:0] _783;
  wire [63:0] _782;
  wire [63:0] _781;
  wire [63:0] _780;
  wire [63:0] _779;
  wire [63:0] _778;
  wire [63:0] _777;
  wire [63:0] _776;
  wire [63:0] _775;
  wire [31:0] _774;
  wire [63:0] _773;
  wire [63:0] _772;
  wire [63:0] _771;
  wire [63:0] _770;
  wire [63:0] _769;
  wire [31:0] _768;
  wire [63:0] _767;
  wire [63:0] _766;
  wire [63:0] _765;
  wire [63:0] _764;
  wire [63:0] _763;
  wire [63:0] _762;
  wire [63:0] _761;
  wire [63:0] _760;
  wire [63:0] _759;
  wire [31:0] _758;
  wire [63:0] _757;
  wire [63:0] _756;
  wire [63:0] _755;
  wire [63:0] _754;
  wire [63:0] _753;
  wire [31:0] _752;
  wire [63:0] _751;
  wire [63:0] _750;
  wire [63:0] _749;
  wire [63:0] _748;
  wire [63:0] _747;
  wire [63:0] _746;
  wire [63:0] _745;
  wire [63:0] _744;
  wire [63:0] _743;
  wire [63:0] _742;
  wire [63:0] _741;
  wire [31:0] _740;
  wire [63:0] _739;
  wire [63:0] _738;
  wire [63:0] _737;
  wire [63:0] _736;
  wire [63:0] _735;
  wire [31:0] _734;
  wire [63:0] _733;
  wire [63:0] _732;
  wire [63:0] _731;
  wire [63:0] _730;
  wire [63:0] _729;
  wire [63:0] _728;
  wire [63:0] _727;
  wire [63:0] _726;
  wire [63:0] _725;
  wire [31:0] _724;
  wire [63:0] _723;
  wire [63:0] _722;
  wire [63:0] _721;
  wire [63:0] _720;
  wire [63:0] _719;
  wire [31:0] _718;
  wire [63:0] _717;
  wire [63:0] _716;
  wire [63:0] _715;
  wire [63:0] _714;
  wire [31:0] _713;
  wire [63:0] _712;
  wire [63:0] _711;
  wire [63:0] _710;
  wire [0:0] ifout752;
  wire [63:0] _709;
  wire [63:0] _708;
  wire [63:0] _707;
  wire [63:0] _706;
  wire [63:0] _705;
  wire [63:0] _704;
  wire [31:0] off_2608;
  wire [31:0] idx_2607;
  wire [31:0] idx_sail_2606;
  wire [31:0] _703;
  wire [31:0] _702;
  wire [63:0] _701;
  wire [31:0] _700;
  wire [31:0] ck_idx_2605;
  wire [31:0] _699;
  wire [63:0] _698;
  wire [63:0] _697;
  wire [63:0] _696;
  wire [63:0] _695;
  wire [63:0] _694;
  wire [63:0] _693;
  wire [63:0] _692;
  wire [63:0] _691;
  wire [63:0] _690;
  wire [63:0] _689;
  wire [63:0] _688;
  wire [63:0] _687;
  wire [31:0] _686;
  wire [63:0] _685;
  wire [63:0] _684;
  wire [63:0] _683;
  wire [63:0] _682;
  wire [63:0] _681;
  wire [31:0] _680;
  wire [63:0] _679;
  wire [63:0] _678;
  wire [63:0] _677;
  wire [63:0] _676;
  wire [63:0] _675;
  wire [63:0] _674;
  wire [63:0] _673;
  wire [63:0] _672;
  wire [63:0] _671;
  wire [31:0] _670;
  wire [63:0] _669;
  wire [63:0] _668;
  wire [63:0] _667;
  wire [63:0] _666;
  wire [63:0] _665;
  wire [31:0] _664;
  wire [63:0] _663;
  wire [63:0] _662;
  wire [63:0] _661;
  wire [63:0] _660;
  wire [63:0] _659;
  wire [63:0] _658;
  wire [63:0] _657;
  wire [63:0] _656;
  wire [63:0] _655;
  wire [63:0] _654;
  wire [63:0] _653;
  wire [31:0] _652;
  wire [63:0] _651;
  wire [63:0] _650;
  wire [63:0] _649;
  wire [63:0] _648;
  wire [63:0] _647;
  wire [31:0] _646;
  wire [63:0] _645;
  wire [63:0] _644;
  wire [63:0] _643;
  wire [63:0] _642;
  wire [63:0] _641;
  wire [63:0] _640;
  wire [63:0] _639;
  wire [63:0] _638;
  wire [63:0] _637;
  wire [31:0] _636;
  wire [63:0] _635;
  wire [63:0] _634;
  wire [63:0] _633;
  wire [63:0] _632;
  wire [63:0] _631;
  wire [31:0] _630;
  wire [63:0] _629;
  wire [63:0] _628;
  wire [63:0] _627;
  wire [63:0] _626;
  wire [31:0] _625;
  wire [63:0] _624;
  wire [63:0] _623;
  wire [63:0] _622;
  wire [0:0] ifout659;
  wire [63:0] _621;
  wire [63:0] _620;
  wire [63:0] _619;
  wire [63:0] _618;
  wire [63:0] _617;
  wire [63:0] _616;
  wire [31:0] off_2598;
  wire [31:0] idx_2597;
  wire [31:0] idx_sail_2596;
  wire [31:0] _615;
  wire [63:0] _614;
  wire [31:0] _613;
  wire [31:0] ck_idx_2594;
  wire [31:0] _612;
  wire [63:0] _611;
  wire [63:0] _610;
  wire [63:0] _609;
  wire [63:0] _608;
  wire [63:0] _607;
  wire [63:0] _606;
  wire [63:0] _605;
  wire [63:0] _604;
  wire [63:0] _603;
  wire [63:0] _602;
  wire [63:0] _601;
  wire [63:0] _600;
  wire [31:0] _599;
  wire [63:0] _598;
  wire [63:0] _597;
  wire [63:0] _596;
  wire [63:0] _595;
  wire [63:0] _594;
  wire [31:0] _593;
  wire [63:0] _592;
  wire [63:0] _591;
  wire [63:0] _590;
  wire [63:0] _589;
  wire [63:0] _588;
  wire [63:0] _587;
  wire [63:0] _586;
  wire [63:0] _585;
  wire [63:0] _584;
  wire [31:0] _583;
  wire [63:0] _582;
  wire [63:0] _581;
  wire [63:0] _580;
  wire [63:0] _579;
  wire [63:0] _578;
  wire [31:0] _577;
  wire [63:0] _576;
  wire [63:0] _575;
  wire [63:0] _574;
  wire [63:0] _573;
  wire [63:0] _572;
  wire [63:0] _571;
  wire [63:0] _570;
  wire [63:0] _569;
  wire [63:0] _568;
  wire [63:0] _567;
  wire [63:0] _566;
  wire [31:0] _565;
  wire [63:0] _564;
  wire [63:0] _563;
  wire [63:0] _562;
  wire [63:0] _561;
  wire [63:0] _560;
  wire [31:0] _559;
  wire [63:0] _558;
  wire [63:0] _557;
  wire [63:0] _556;
  wire [63:0] _555;
  wire [63:0] _554;
  wire [63:0] _553;
  wire [63:0] _552;
  wire [63:0] _551;
  wire [63:0] _550;
  wire [31:0] _549;
  wire [63:0] _548;
  wire [63:0] _547;
  wire [63:0] _546;
  wire [63:0] _545;
  wire [63:0] _544;
  wire [31:0] _543;
  wire [63:0] _542;
  wire [63:0] _541;
  wire [63:0] _540;
  wire [63:0] _539;
  wire [31:0] _538;
  wire [63:0] _537;
  wire [63:0] _536;
  wire [63:0] _535;
  wire [0:0] ifout567;
  wire [63:0] _534;
  wire [63:0] _533;
  wire [63:0] _532;
  wire [63:0] _531;
  wire [63:0] _530;
  wire [63:0] _529;
  wire [31:0] off_2587;
  wire [31:0] idx_2586;
  wire [31:0] idx_sail_2585;
  wire [31:0] _528;
  wire [31:0] _527;
  wire [31:0] _526;
  wire [31:0] ck_idx_2584;
  wire [31:0] _525;
  wire [63:0] _524;
  wire [63:0] _523;
  wire [63:0] _522;
  wire [63:0] _521;
  wire [63:0] _520;
  wire [63:0] _519;
  wire [63:0] _518;
  wire [63:0] _517;
  wire [63:0] _516;
  wire [63:0] _515;
  wire [63:0] _514;
  wire [63:0] _513;
  wire [31:0] _512;
  wire [63:0] _511;
  wire [63:0] _510;
  wire [63:0] _509;
  wire [63:0] _508;
  wire [63:0] _507;
  wire [31:0] _506;
  wire [63:0] _505;
  wire [63:0] _504;
  wire [63:0] _503;
  wire [63:0] _502;
  wire [63:0] _501;
  wire [63:0] _500;
  wire [63:0] _499;
  wire [63:0] _498;
  wire [63:0] _497;
  wire [31:0] _496;
  wire [63:0] _495;
  wire [63:0] _494;
  wire [63:0] _493;
  wire [63:0] _492;
  wire [63:0] _491;
  wire [31:0] _490;
  wire [63:0] _489;
  wire [63:0] _488;
  wire [63:0] _487;
  wire [63:0] _486;
  wire [63:0] _485;
  wire [63:0] _484;
  wire [63:0] _483;
  wire [63:0] _482;
  wire [63:0] _481;
  wire [63:0] _480;
  wire [63:0] _479;
  wire [31:0] _478;
  wire [63:0] _477;
  wire [63:0] _476;
  wire [63:0] _475;
  wire [63:0] _474;
  wire [63:0] _473;
  wire [31:0] _472;
  wire [63:0] _471;
  wire [63:0] _470;
  wire [63:0] _469;
  wire [63:0] _468;
  wire [63:0] _467;
  wire [63:0] _466;
  wire [63:0] _465;
  wire [63:0] _464;
  wire [63:0] _463;
  wire [31:0] _462;
  wire [63:0] _461;
  wire [63:0] _460;
  wire [63:0] _459;
  wire [63:0] _458;
  wire [63:0] _457;
  wire [31:0] _456;
  wire [63:0] _455;
  wire [63:0] _454;
  wire [63:0] _453;
  wire [63:0] _452;
  wire [31:0] _451;
  wire [63:0] _450;
  wire [63:0] _449;
  wire [63:0] _448;
  wire [0:0] ifout475;
  wire [63:0] _447;
  wire [63:0] _446;
  wire [63:0] _445;
  wire [63:0] _444;
  wire [63:0] _443;
  wire [63:0] _442;
  wire [31:0] off_2577;
  wire [31:0] idx_2576;
  wire [31:0] idx_sail_2575;
  wire [31:0] _441;
  wire [31:0] _440;
  wire [63:0] _439;
  wire [31:0] _438;
  wire [31:0] ck_idx_2574;
  wire [31:0] _437;
  wire [63:0] _436;
  wire [63:0] _435;
  wire [63:0] _434;
  wire [63:0] _433;
  wire [63:0] _432;
  wire [63:0] _431;
  wire [63:0] _430;
  wire [63:0] _429;
  wire [63:0] _428;
  wire [63:0] _427;
  wire [63:0] _426;
  wire [63:0] _425;
  wire [31:0] _424;
  wire [63:0] _423;
  wire [63:0] _422;
  wire [63:0] _421;
  wire [63:0] _420;
  wire [63:0] _419;
  wire [31:0] _418;
  wire [63:0] _417;
  wire [63:0] _416;
  wire [63:0] _415;
  wire [63:0] _414;
  wire [63:0] _413;
  wire [63:0] _412;
  wire [63:0] _411;
  wire [63:0] _410;
  wire [63:0] _409;
  wire [31:0] _408;
  wire [63:0] _407;
  wire [63:0] _406;
  wire [63:0] _405;
  wire [63:0] _404;
  wire [63:0] _403;
  wire [31:0] _402;
  wire [63:0] _401;
  wire [63:0] _400;
  wire [63:0] _399;
  wire [63:0] _398;
  wire [63:0] _397;
  wire [63:0] _396;
  wire [63:0] _395;
  wire [63:0] _394;
  wire [63:0] _393;
  wire [63:0] _392;
  wire [63:0] _391;
  wire [31:0] _390;
  wire [63:0] _389;
  wire [63:0] _388;
  wire [63:0] _387;
  wire [63:0] _386;
  wire [63:0] _385;
  wire [31:0] _384;
  wire [63:0] _383;
  wire [63:0] _382;
  wire [63:0] _381;
  wire [63:0] _380;
  wire [63:0] _379;
  wire [63:0] _378;
  wire [63:0] _377;
  wire [63:0] _376;
  wire [63:0] _375;
  wire [31:0] _374;
  wire [63:0] _373;
  wire [63:0] _372;
  wire [63:0] _371;
  wire [63:0] _370;
  wire [63:0] _369;
  wire [31:0] _368;
  wire [63:0] _367;
  wire [63:0] _366;
  wire [63:0] _365;
  wire [63:0] _364;
  wire [31:0] _363;
  wire [63:0] _362;
  wire [63:0] _361;
  wire [63:0] _360;
  wire [0:0] ifout382;
  wire [63:0] _359;
  wire [63:0] _358;
  wire [63:0] _357;
  wire [63:0] _356;
  wire [63:0] _355;
  wire [63:0] _354;
  wire [31:0] off_2567;
  wire [31:0] idx_2566;
  wire [31:0] idx_sail_2565;
  wire [31:0] _353;
  wire [31:0] _352;
  wire [63:0] _351;
  wire [31:0] _350;
  wire [31:0] ck_idx_2564;
  wire [31:0] _349;
  wire [63:0] _348;
  wire [63:0] _347;
  wire [63:0] _346;
  wire [63:0] _345;
  wire [63:0] _344;
  wire [63:0] _343;
  wire [63:0] _342;
  wire [63:0] _341;
  wire [63:0] _340;
  wire [63:0] _339;
  wire [63:0] _338;
  wire [63:0] _337;
  wire [31:0] _336;
  wire [63:0] _335;
  wire [63:0] _334;
  wire [63:0] _333;
  wire [63:0] _332;
  wire [63:0] _331;
  wire [31:0] _330;
  wire [63:0] _329;
  wire [63:0] _328;
  wire [63:0] _327;
  wire [63:0] _326;
  wire [63:0] _325;
  wire [63:0] _324;
  wire [63:0] _323;
  wire [63:0] _322;
  wire [63:0] _321;
  wire [31:0] _320;
  wire [63:0] _319;
  wire [63:0] _318;
  wire [63:0] _317;
  wire [63:0] _316;
  wire [63:0] _315;
  wire [31:0] _314;
  wire [63:0] _313;
  wire [63:0] _312;
  wire [63:0] _311;
  wire [63:0] _310;
  wire [63:0] _309;
  wire [63:0] _308;
  wire [63:0] _307;
  wire [63:0] _306;
  wire [63:0] _305;
  wire [63:0] _304;
  wire [63:0] _303;
  wire [31:0] _302;
  wire [63:0] _301;
  wire [63:0] _300;
  wire [63:0] _299;
  wire [63:0] _298;
  wire [63:0] _297;
  wire [31:0] _296;
  wire [63:0] _295;
  wire [63:0] _294;
  wire [63:0] _293;
  wire [63:0] _292;
  wire [63:0] _291;
  wire [63:0] _290;
  wire [63:0] _289;
  wire [63:0] _288;
  wire [63:0] _287;
  wire [31:0] _286;
  wire [63:0] _285;
  wire [63:0] _284;
  wire [63:0] _283;
  wire [63:0] _282;
  wire [63:0] _281;
  wire [31:0] _280;
  wire [63:0] _279;
  wire [63:0] _278;
  wire [63:0] _277;
  wire [63:0] _276;
  wire [31:0] _275;
  wire [63:0] _274;
  wire [63:0] _273;
  wire [63:0] _272;
  wire [0:0] ifout289;
  wire [63:0] _271;
  wire [63:0] _270;
  wire [63:0] _269;
  wire [63:0] _268;
  wire [63:0] _267;
  wire [63:0] _266;
  wire [31:0] off_2557;
  wire [31:0] idx_2556;
  wire [31:0] idx_sail_2555;
  wire [31:0] _265;
  wire [31:0] _264;
  wire [63:0] _263;
  wire [31:0] _262;
  wire [31:0] ck_idx_2554;
  wire [31:0] _261;
  wire [63:0] _260;
  wire [63:0] _259;
  wire [63:0] _258;
  wire [63:0] _257;
  wire [63:0] _256;
  wire [63:0] _255;
  wire [63:0] _254;
  wire [63:0] _253;
  wire [63:0] _252;
  wire [63:0] _251;
  wire [63:0] _250;
  wire [63:0] _249;
  wire [31:0] _248;
  wire [63:0] _247;
  wire [63:0] _246;
  wire [63:0] _245;
  wire [63:0] _244;
  wire [63:0] _243;
  wire [31:0] _242;
  wire [63:0] _241;
  wire [63:0] _240;
  wire [63:0] _239;
  wire [63:0] _238;
  wire [63:0] _237;
  wire [63:0] _236;
  wire [63:0] _235;
  wire [63:0] _234;
  wire [63:0] _233;
  wire [31:0] _232;
  wire [63:0] _231;
  wire [63:0] _230;
  wire [63:0] _229;
  wire [63:0] _228;
  wire [63:0] _227;
  wire [31:0] _226;
  wire [63:0] _225;
  wire [63:0] _224;
  wire [63:0] _223;
  wire [63:0] _222;
  wire [63:0] _221;
  wire [63:0] _220;
  wire [63:0] _219;
  wire [63:0] _218;
  wire [63:0] _217;
  wire [63:0] _216;
  wire [63:0] _215;
  wire [31:0] _214;
  wire [63:0] _213;
  wire [63:0] _212;
  wire [63:0] _211;
  wire [63:0] _210;
  wire [63:0] _209;
  wire [31:0] _208;
  wire [63:0] _207;
  wire [63:0] _206;
  wire [63:0] _205;
  wire [63:0] _204;
  wire [63:0] _203;
  wire [63:0] _202;
  wire [63:0] _201;
  wire [63:0] _200;
  wire [63:0] _199;
  wire [31:0] _198;
  wire [63:0] _197;
  wire [63:0] _196;
  wire [63:0] _195;
  wire [63:0] _194;
  wire [63:0] _193;
  wire [31:0] _192;
  wire [63:0] _191;
  wire [63:0] _190;
  wire [63:0] _189;
  wire [63:0] _188;
  wire [31:0] _187;
  wire [63:0] _186;
  wire [63:0] _185;
  wire [63:0] _184;
  wire [0:0] ifout196;
  wire [63:0] _183;
  wire [63:0] _182;
  wire [63:0] _181;
  wire [63:0] _180;
  wire [63:0] _179;
  wire [63:0] _178;
  wire [31:0] off_2547;
  wire [31:0] idx_2546;
  wire [31:0] idx_sail_2545;
  wire [31:0] _177;
  wire [31:0] _176;
  wire [63:0] _175;
  wire [31:0] _174;
  wire [31:0] ck_idx_2544;
  wire [31:0] _173;
  wire [63:0] _172;
  wire [63:0] _171;
  wire [63:0] _170;
  wire [63:0] _169;
  wire [63:0] _168;
  wire [63:0] _167;
  wire [63:0] _166;
  wire [63:0] _165;
  wire [63:0] _164;
  wire [63:0] _163;
  wire [63:0] _162;
  wire [63:0] _161;
  wire [31:0] _160;
  wire [63:0] _159;
  wire [63:0] _158;
  wire [63:0] _157;
  wire [63:0] _156;
  wire [63:0] _155;
  wire [31:0] _154;
  wire [63:0] _153;
  wire [63:0] _152;
  wire [63:0] _151;
  wire [63:0] _150;
  wire [63:0] _149;
  wire [63:0] _148;
  wire [63:0] _147;
  wire [63:0] _146;
  wire [63:0] _145;
  wire [31:0] _144;
  wire [63:0] _143;
  wire [63:0] _142;
  wire [63:0] _141;
  wire [63:0] _140;
  wire [63:0] _139;
  wire [31:0] _138;
  wire [63:0] _137;
  wire [63:0] _136;
  wire [63:0] _135;
  wire [63:0] _134;
  wire [63:0] _133;
  wire [63:0] _132;
  wire [63:0] _131;
  wire [63:0] _130;
  wire [63:0] _129;
  wire [63:0] _128;
  wire [63:0] _127;
  wire [31:0] _126;
  wire [63:0] _125;
  wire [63:0] _124;
  wire [63:0] _123;
  wire [63:0] _122;
  wire [63:0] _121;
  wire [31:0] _120;
  wire [63:0] _119;
  wire [63:0] _118;
  wire [63:0] _117;
  wire [63:0] _116;
  wire [63:0] _115;
  wire [63:0] _114;
  wire [63:0] _113;
  wire [63:0] _112;
  wire [63:0] _111;
  wire [31:0] _110;
  wire [63:0] _109;
  wire [63:0] _108;
  wire [63:0] _107;
  wire [63:0] _106;
  wire [63:0] _105;
  wire [31:0] _104;
  wire [63:0] _103;
  wire [63:0] _102;
  wire [63:0] _101;
  wire [63:0] _100;
  wire [31:0] _99;
  wire [63:0] _98;
  wire [63:0] _97;
  wire [63:0] _96;
  wire [0:0] ifout103;
  wire [63:0] _95;
  wire [63:0] _94;
  wire [63:0] _93;
  wire [63:0] _92;
  wire [63:0] _91;
  wire [63:0] _90;
  wire [31:0] off_2537;
  wire [31:0] idx_2536;
  wire [31:0] idx_sail_2535;
  wire [31:0] _89;
  wire [31:0] _88;
  wire [63:0] _87;
  wire [31:0] _86;
  wire [31:0] ck_idx_2534;
  wire [31:0] _85;
  wire [63:0] _84;
  wire [63:0] _83;
  wire [63:0] _82;
  wire [63:0] _81;
  wire [63:0] _80;
  wire [63:0] _79;
  wire [63:0] _78;
  wire [63:0] _77;
  wire [63:0] _76;
  wire [63:0] _75;
  wire [63:0] _74;
  wire [63:0] _73;
  wire [31:0] _72;
  wire [63:0] _71;
  wire [63:0] _70;
  wire [63:0] _69;
  wire [63:0] _68;
  wire [63:0] _67;
  wire [31:0] _66;
  wire [63:0] _65;
  wire [63:0] _64;
  wire [63:0] _63;
  wire [63:0] _62;
  wire [63:0] _61;
  wire [63:0] _60;
  wire [63:0] _59;
  wire [63:0] _58;
  wire [63:0] _57;
  wire [31:0] _56;
  wire [63:0] _55;
  wire [63:0] _54;
  wire [63:0] _53;
  wire [63:0] _52;
  wire [63:0] _51;
  wire [31:0] _50;
  wire [63:0] _49;
  wire [63:0] _48;
  wire [63:0] _47;
  wire [63:0] _46;
  wire [63:0] _45;
  wire [63:0] _44;
  wire [63:0] _43;
  wire [63:0] _42;
  wire [63:0] _41;
  wire [63:0] _40;
  wire [63:0] _39;
  wire [31:0] _38;
  wire [63:0] _37;
  wire [63:0] _36;
  wire [63:0] _35;
  wire [63:0] _34;
  wire [63:0] _33;
  wire [31:0] _32;
  wire [63:0] _31;
  wire [63:0] _30;
  wire [63:0] _29;
  wire [63:0] _28;
  wire [63:0] _27;
  wire [63:0] _26;
  wire [63:0] _25;
  wire [63:0] _24;
  wire [63:0] _23;
  wire [31:0] _22;
  wire [63:0] _21;
  wire [63:0] _20;
  wire [63:0] _19;
  wire [63:0] _18;
  wire [63:0] _17;
  wire [31:0] _16;
  wire [63:0] _15;
  wire [63:0] _14;
  wire [63:0] _13;
  wire [63:0] _12;
  wire [31:0] _11;
  wire [63:0] _10;
  wire [63:0] _9;
  wire [63:0] _8;
  wire [0:0] ifout10;
  wire [63:0] _7;
  wire [63:0] _6;
  wire [63:0] _5;
  wire [63:0] _4;
  wire [63:0] _3;
  wire [63:0] _2;
  wire [31:0] off_2525;
  wire [31:0] idx_2524;
  wire [31:0] idx_sail_2523;
  wire [63:0] _1;
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op0 (.out1(_1), .in1(ip1_2522_D), .in2(6 'd 48));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1 (.out1(idx_sail_2523), .in1(_1));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(3), .BITSIZE_out1(32), .PRECISION(32)) op2 (.out1(idx_2524), .in1(idx_sail_2523), .in2(3 'd 6));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2668 (.out1(R2669), .clock(clock), .in1(idx_sail_2523));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2671 (.out1(R2672), .clock(clock), .in1(idx_2524));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op4 (.out1(_2), .in1(R2672));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op5 (.out1(_3), .in1(_2), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2669 (.out1(R2670), .clock(clock), .in1(R2669));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2672 (.out1(R2673), .clock(clock), .in1(R2672));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2877 (.out1(R2878), .clock(clock), .in1(_3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op6 (.out1(_4), .in1(c16_bitmap_2526_D), .in2(R2878));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2670 (.out1(R2671), .clock(clock), .in1(R2670));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2673 (.out1(R2674), .clock(clock), .in1(R2673));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2878 (.out1(R2879), .clock(clock), .in1(_4));
  SRAM op7 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_5),.ADR(R2879));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op3 (.out1(off_2525), .in1(R2671), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op8 (.out1(_6), .in1(64 'd 9223372036854775808), .in2(off_2525));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2674 (.out1(R2675), .clock(clock), .in1(R2674));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op2879 (.out1(R2880), .clock(clock), .in1(_5));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2880 (.out1(R2881), .clock(clock), .in1(off_2525));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3082 (.out1(R3083), .clock(clock), .in1(_6));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op9 (.out1(_7), .in1(R2880), .in2(R3083));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op10 (.out1(ifout10), .in1(_7), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op71 (.out1(_68), .in1(R2675));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op72 (.out1(_69), .in1(_68), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2675 (.out1(R2676), .clock(clock), .in1(R2675));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2881 (.out1(R2882), .clock(clock), .in1(R2881));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3083 (.out1(R3084), .clock(clock), .in1(ifout10));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3291 (.out1(R3292), .clock(clock), .in1(_69));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op65 (.out1(_62), .in1(R2676));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op55 (.out1(_52), .in1(R2676));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op49 (.out1(_46), .in1(R2676));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op37 (.out1(_34), .in1(R2676));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op31 (.out1(_28), .in1(R2676));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op21 (.out1(_18), .in1(R2676));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op66 (.out1(_63), .in1(_62), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op56 (.out1(_53), .in1(_52), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op50 (.out1(_47), .in1(_46), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op38 (.out1(_35), .in1(_34), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op32 (.out1(_29), .in1(_28), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op22 (.out1(_19), .in1(_18), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op73 (.out1(_70), .in1(c16_bitmap_2526_D), .in2(R3292));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2676 (.out1(R2677), .clock(clock), .in1(R2676));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2882 (.out1(R2883), .clock(clock), .in1(R2882));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3084 (.out1(R3085), .clock(clock), .in1(R3084));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3292 (.out1(R3293), .clock(clock), .in1(_63));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3293 (.out1(R3294), .clock(clock), .in1(_53));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3294 (.out1(R3295), .clock(clock), .in1(_47));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3295 (.out1(R3296), .clock(clock), .in1(_35));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3296 (.out1(R3297), .clock(clock), .in1(_29));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3297 (.out1(R3298), .clock(clock), .in1(_19));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3298 (.out1(R3299), .clock(clock), .in1(_70));
  SRAM op74 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_71),.ADR(R3299));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op15 (.out1(_12), .in1(R2677));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op16 (.out1(_13), .in1(_12), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op67 (.out1(_64), .in1(c16_bitmap_2526_D), .in2(R3293));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op57 (.out1(_54), .in1(c16_bitmap_2526_D), .in2(R3294));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op51 (.out1(_48), .in1(c16_bitmap_2526_D), .in2(R3295));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op39 (.out1(_36), .in1(c16_bitmap_2526_D), .in2(R3296));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op33 (.out1(_30), .in1(c16_bitmap_2526_D), .in2(R3297));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op23 (.out1(_20), .in1(c16_bitmap_2526_D), .in2(R3298));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2677 (.out1(R2678), .clock(clock), .in1(R2677));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2883 (.out1(R2884), .clock(clock), .in1(R2883));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3085 (.out1(R3086), .clock(clock), .in1(R3085));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3299 (.out1(R3300), .clock(clock), .in1(_71));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3300 (.out1(R3301), .clock(clock), .in1(_13));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3301 (.out1(R3302), .clock(clock), .in1(_64));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3302 (.out1(R3303), .clock(clock), .in1(_54));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3303 (.out1(R3304), .clock(clock), .in1(_48));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3304 (.out1(R3305), .clock(clock), .in1(_36));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3305 (.out1(R3306), .clock(clock), .in1(_30));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3306 (.out1(R3307), .clock(clock), .in1(_20));
  SRAM op68 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_65),.ADR(R3302));
  SRAM op58 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_55),.ADR(R3303));
  SRAM op52 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_49),.ADR(R3304));
  SRAM op40 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_37),.ADR(R3305));
  SRAM op34 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_31),.ADR(R3306));
  SRAM op24 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_21),.ADR(R3307));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op75 (.out1(_72), .in1(7 'd 64), .in2(R2884));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op17 (.out1(_14), .in1(c16_bitmap_2526_D), .in2(R3301));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op76 (.out1(_73), .in1(R3300), .in2(_72));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op69 (.out1(_66), .in1(7 'd 64), .in2(R2884));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op59 (.out1(_56), .in1(7 'd 64), .in2(R2884));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op41 (.out1(_38), .in1(7 'd 64), .in2(R2884));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2678 (.out1(R2679), .clock(clock), .in1(R2678));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2884 (.out1(R2885), .clock(clock), .in1(R2884));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3086 (.out1(R3087), .clock(clock), .in1(R3086));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3307 (.out1(R3308), .clock(clock), .in1(_65));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3308 (.out1(R3309), .clock(clock), .in1(_55));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3309 (.out1(R3310), .clock(clock), .in1(_49));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3310 (.out1(R3311), .clock(clock), .in1(_37));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3311 (.out1(R3312), .clock(clock), .in1(_31));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3312 (.out1(R3313), .clock(clock), .in1(_21));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3313 (.out1(R3314), .clock(clock), .in1(_14));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3314 (.out1(R3315), .clock(clock), .in1(_73));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3315 (.out1(R3316), .clock(clock), .in1(_66));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3316 (.out1(R3317), .clock(clock), .in1(_56));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3317 (.out1(R3318), .clock(clock), .in1(_38));
  SRAM op18 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_15),.ADR(R3314));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op77 (.out1(_74), .in1(R3315), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op70 (.out1(_67), .in1(R3308), .in2(R3316));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op60 (.out1(_57), .in1(R3309), .in2(R3317));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op53 (.out1(_50), .in1(7 'd 64), .in2(R2885));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op42 (.out1(_39), .in1(R3311), .in2(R3318));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op35 (.out1(_32), .in1(7 'd 64), .in2(R2885));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op25 (.out1(_22), .in1(7 'd 64), .in2(R2885));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op78 (.out1(_75), .in1(_74), .in2(63 'd 6148914691236517205));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op79 (.out1(_76), .in1(_67), .in2(_75));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op61 (.out1(_58), .in1(_57), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op54 (.out1(_51), .in1(R3310), .in2(_50));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op43 (.out1(_40), .in1(_39), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op36 (.out1(_33), .in1(R3312), .in2(_32));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op26 (.out1(_23), .in1(R3313), .in2(_22));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op19 (.out1(_16), .in1(7 'd 64), .in2(R2885));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2679 (.out1(R2680), .clock(clock), .in1(R2679));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2885 (.out1(R2886), .clock(clock), .in1(R2885));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3087 (.out1(R3088), .clock(clock), .in1(R3087));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3318 (.out1(R3319), .clock(clock), .in1(_15));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3319 (.out1(R3320), .clock(clock), .in1(_76));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3320 (.out1(R3321), .clock(clock), .in1(_58));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3321 (.out1(R3322), .clock(clock), .in1(_51));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3322 (.out1(R3323), .clock(clock), .in1(_40));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3323 (.out1(R3324), .clock(clock), .in1(_33));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3324 (.out1(R3325), .clock(clock), .in1(_23));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3325 (.out1(R3326), .clock(clock), .in1(_16));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op11 (.out1(_8), .in1(R2680));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op62 (.out1(_59), .in1(R3321), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op80 (.out1(_77), .in1(R3320), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op63 (.out1(_60), .in1(R3322), .in2(_59));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op44 (.out1(_41), .in1(R3323), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op27 (.out1(_24), .in1(R3325), .in2(1 'd 1));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op45 (.out1(_42), .in1(R3324), .in2(_41));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op20 (.out1(_17), .in1(R3319), .in2(R3326));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op12 (.out1(_9), .in1(_8), .in2(2 'd 2));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op81 (.out1(_78), .in1(_77), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op64 (.out1(_61), .in1(_60), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op28 (.out1(_25), .in1(_24), .in2(63 'd 6148914691236517205));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op82 (.out1(_79), .in1(_61), .in2(_78));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op46 (.out1(_43), .in1(_42), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op29 (.out1(_26), .in1(_17), .in2(_25));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2680 (.out1(R2681), .clock(clock), .in1(R2680));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2886 (.out1(R2887), .clock(clock), .in1(R2886));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3088 (.out1(R3089), .clock(clock), .in1(R3088));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3326 (.out1(R3327), .clock(clock), .in1(_9));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3327 (.out1(R3328), .clock(clock), .in1(_79));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3328 (.out1(R3329), .clock(clock), .in1(_43));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3329 (.out1(R3330), .clock(clock), .in1(_26));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op47 (.out1(_44), .in1(R3329), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op30 (.out1(_27), .in1(R3330), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op83 (.out1(_80), .in1(R3328), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op48 (.out1(_45), .in1(_27), .in2(_44));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op13 (.out1(_10), .in1(c16_popcnt_2533_D), .in2(R3327));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op84 (.out1(_81), .in1(_45), .in2(_80));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op85 (.out1(_82), .in1(_81), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2681 (.out1(R2682), .clock(clock), .in1(R2681));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2887 (.out1(R2888), .clock(clock), .in1(R2887));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3089 (.out1(R3090), .clock(clock), .in1(R3089));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3330 (.out1(R3331), .clock(clock), .in1(_10));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3331 (.out1(R3332), .clock(clock), .in1(_82));
  SRAM op14 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_11),.ADR(R3331));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op86 (.out1(_83), .in1(R3332), .in2(57 'd 72340172838076673));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2682 (.out1(R2683), .clock(clock), .in1(R2682));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2888 (.out1(R2889), .clock(clock), .in1(R2888));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3090 (.out1(R3091), .clock(clock), .in1(R3090));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3332 (.out1(R3333), .clock(clock), .in1(_11));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3333 (.out1(R3334), .clock(clock), .in1(_83));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op87 (.out1(_84), .in1(R3334), .in2(6 'd 56));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op88 (.out1(_85), .in1(_84));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op89 (.out1(ck_idx_2534), .in1(R3333), .in2(_85));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2683 (.out1(R2684), .clock(clock), .in1(R2683));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2889 (.out1(R2890), .clock(clock), .in1(R2889));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3091 (.out1(R3092), .clock(clock), .in1(R3091));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3334 (.out1(R3335), .clock(clock), .in1(ck_idx_2534));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(4), .BITSIZE_out1(32), .PRECISION(32)) op90 (.out1(_86), .in1(R3335), .in2(4 'd 8));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op91 (.out1(_87), .in1(ip1_2522_D), .in2(6 'd 40));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2684 (.out1(R2685), .clock(clock), .in1(R2684));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2890 (.out1(R2891), .clock(clock), .in1(R2890));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3092 (.out1(R3093), .clock(clock), .in1(R3092));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3335 (.out1(R3336), .clock(clock), .in1(_86));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3336 (.out1(R3337), .clock(clock), .in1(_87));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op92 (.out1(_88), .in1(R3337));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(8), .BITSIZE_out1(32)) op93 (.out1(_89), .in1(_88), .in2(8 'd 255));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op94 (.out1(idx_sail_2535), .in1(R3336), .in2(_89));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(3), .BITSIZE_out1(32), .PRECISION(32)) op95 (.out1(idx_2536), .in1(idx_sail_2535), .in2(3 'd 6));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2685 (.out1(R2686), .clock(clock), .in1(R2685));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2891 (.out1(R2892), .clock(clock), .in1(R2891));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3093 (.out1(R3094), .clock(clock), .in1(R3093));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3337 (.out1(R3338), .clock(clock), .in1(idx_sail_2535));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3340 (.out1(R3341), .clock(clock), .in1(idx_2536));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op97 (.out1(_90), .in1(R3341));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op98 (.out1(_91), .in1(_90), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2686 (.out1(R2687), .clock(clock), .in1(R2686));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2892 (.out1(R2893), .clock(clock), .in1(R2892));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3094 (.out1(R3095), .clock(clock), .in1(R3094));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3338 (.out1(R3339), .clock(clock), .in1(R3338));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3341 (.out1(R3342), .clock(clock), .in1(R3341));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3532 (.out1(R3533), .clock(clock), .in1(_91));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op99 (.out1(_92), .in1(c24_bitmap_2538_D), .in2(R3533));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2687 (.out1(R2688), .clock(clock), .in1(R2687));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2893 (.out1(R2894), .clock(clock), .in1(R2893));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3095 (.out1(R3096), .clock(clock), .in1(R3095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3339 (.out1(R3340), .clock(clock), .in1(R3339));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3342 (.out1(R3343), .clock(clock), .in1(R3342));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3533 (.out1(R3534), .clock(clock), .in1(_92));
  SRAM op100 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_93),.ADR(R3534));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op96 (.out1(off_2537), .in1(R3340), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op101 (.out1(_94), .in1(64 'd 9223372036854775808), .in2(off_2537));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2688 (.out1(R2689), .clock(clock), .in1(R2688));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2894 (.out1(R2895), .clock(clock), .in1(R2894));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3096 (.out1(R3097), .clock(clock), .in1(R3096));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3343 (.out1(R3344), .clock(clock), .in1(R3343));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3534 (.out1(R3535), .clock(clock), .in1(_93));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3535 (.out1(R3536), .clock(clock), .in1(off_2537));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3723 (.out1(R3724), .clock(clock), .in1(_94));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op102 (.out1(_95), .in1(R3535), .in2(R3724));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op103 (.out1(ifout103), .in1(_95), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op164 (.out1(_156), .in1(R3344));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op165 (.out1(_157), .in1(_156), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2689 (.out1(R2690), .clock(clock), .in1(R2689));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2895 (.out1(R2896), .clock(clock), .in1(R2895));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3097 (.out1(R3098), .clock(clock), .in1(R3097));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3344 (.out1(R3345), .clock(clock), .in1(R3344));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3536 (.out1(R3537), .clock(clock), .in1(R3536));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3724 (.out1(R3725), .clock(clock), .in1(ifout103));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3918 (.out1(R3919), .clock(clock), .in1(_157));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op158 (.out1(_150), .in1(R3345));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op148 (.out1(_140), .in1(R3345));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op142 (.out1(_134), .in1(R3345));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op130 (.out1(_122), .in1(R3345));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op124 (.out1(_116), .in1(R3345));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op114 (.out1(_106), .in1(R3345));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op159 (.out1(_151), .in1(_150), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op149 (.out1(_141), .in1(_140), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op143 (.out1(_135), .in1(_134), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op131 (.out1(_123), .in1(_122), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op125 (.out1(_117), .in1(_116), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op115 (.out1(_107), .in1(_106), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op166 (.out1(_158), .in1(c24_bitmap_2538_D), .in2(R3919));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2690 (.out1(R2691), .clock(clock), .in1(R2690));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2896 (.out1(R2897), .clock(clock), .in1(R2896));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3098 (.out1(R3099), .clock(clock), .in1(R3098));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3345 (.out1(R3346), .clock(clock), .in1(R3345));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3537 (.out1(R3538), .clock(clock), .in1(R3537));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3725 (.out1(R3726), .clock(clock), .in1(R3725));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3919 (.out1(R3920), .clock(clock), .in1(_151));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3920 (.out1(R3921), .clock(clock), .in1(_141));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3921 (.out1(R3922), .clock(clock), .in1(_135));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3922 (.out1(R3923), .clock(clock), .in1(_123));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3923 (.out1(R3924), .clock(clock), .in1(_117));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3924 (.out1(R3925), .clock(clock), .in1(_107));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3925 (.out1(R3926), .clock(clock), .in1(_158));
  SRAM op167 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_159),.ADR(R3926));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op108 (.out1(_100), .in1(R3346));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op109 (.out1(_101), .in1(_100), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op160 (.out1(_152), .in1(c24_bitmap_2538_D), .in2(R3920));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op150 (.out1(_142), .in1(c24_bitmap_2538_D), .in2(R3921));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op144 (.out1(_136), .in1(c24_bitmap_2538_D), .in2(R3922));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op132 (.out1(_124), .in1(c24_bitmap_2538_D), .in2(R3923));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op126 (.out1(_118), .in1(c24_bitmap_2538_D), .in2(R3924));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op116 (.out1(_108), .in1(c24_bitmap_2538_D), .in2(R3925));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2691 (.out1(R2692), .clock(clock), .in1(R2691));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2897 (.out1(R2898), .clock(clock), .in1(R2897));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3099 (.out1(R3100), .clock(clock), .in1(R3099));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3346 (.out1(R3347), .clock(clock), .in1(R3346));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3538 (.out1(R3539), .clock(clock), .in1(R3538));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3726 (.out1(R3727), .clock(clock), .in1(R3726));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3926 (.out1(R3927), .clock(clock), .in1(_159));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3927 (.out1(R3928), .clock(clock), .in1(_101));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3928 (.out1(R3929), .clock(clock), .in1(_152));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3929 (.out1(R3930), .clock(clock), .in1(_142));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3930 (.out1(R3931), .clock(clock), .in1(_136));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3931 (.out1(R3932), .clock(clock), .in1(_124));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3932 (.out1(R3933), .clock(clock), .in1(_118));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3933 (.out1(R3934), .clock(clock), .in1(_108));
  SRAM op161 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_153),.ADR(R3929));
  SRAM op151 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_143),.ADR(R3930));
  SRAM op145 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_137),.ADR(R3931));
  SRAM op133 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_125),.ADR(R3932));
  SRAM op127 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_119),.ADR(R3933));
  SRAM op117 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_109),.ADR(R3934));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op168 (.out1(_160), .in1(7 'd 64), .in2(R3539));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op110 (.out1(_102), .in1(c24_bitmap_2538_D), .in2(R3928));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op169 (.out1(_161), .in1(R3927), .in2(_160));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op162 (.out1(_154), .in1(7 'd 64), .in2(R3539));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op152 (.out1(_144), .in1(7 'd 64), .in2(R3539));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op134 (.out1(_126), .in1(7 'd 64), .in2(R3539));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2692 (.out1(R2693), .clock(clock), .in1(R2692));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2898 (.out1(R2899), .clock(clock), .in1(R2898));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3100 (.out1(R3101), .clock(clock), .in1(R3100));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3347 (.out1(R3348), .clock(clock), .in1(R3347));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3539 (.out1(R3540), .clock(clock), .in1(R3539));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3727 (.out1(R3728), .clock(clock), .in1(R3727));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3934 (.out1(R3935), .clock(clock), .in1(_153));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3935 (.out1(R3936), .clock(clock), .in1(_143));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3936 (.out1(R3937), .clock(clock), .in1(_137));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3937 (.out1(R3938), .clock(clock), .in1(_125));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3938 (.out1(R3939), .clock(clock), .in1(_119));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3939 (.out1(R3940), .clock(clock), .in1(_109));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3940 (.out1(R3941), .clock(clock), .in1(_102));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3941 (.out1(R3942), .clock(clock), .in1(_161));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3942 (.out1(R3943), .clock(clock), .in1(_154));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3943 (.out1(R3944), .clock(clock), .in1(_144));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3944 (.out1(R3945), .clock(clock), .in1(_126));
  SRAM op111 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_103),.ADR(R3941));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op170 (.out1(_162), .in1(R3942), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op163 (.out1(_155), .in1(R3935), .in2(R3943));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op153 (.out1(_145), .in1(R3936), .in2(R3944));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op146 (.out1(_138), .in1(7 'd 64), .in2(R3540));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op135 (.out1(_127), .in1(R3938), .in2(R3945));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op128 (.out1(_120), .in1(7 'd 64), .in2(R3540));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op118 (.out1(_110), .in1(7 'd 64), .in2(R3540));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op171 (.out1(_163), .in1(_162), .in2(63 'd 6148914691236517205));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op172 (.out1(_164), .in1(_155), .in2(_163));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op154 (.out1(_146), .in1(_145), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op147 (.out1(_139), .in1(R3937), .in2(_138));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op136 (.out1(_128), .in1(_127), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op129 (.out1(_121), .in1(R3939), .in2(_120));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op119 (.out1(_111), .in1(R3940), .in2(_110));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op112 (.out1(_104), .in1(7 'd 64), .in2(R3540));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2693 (.out1(R2694), .clock(clock), .in1(R2693));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2899 (.out1(R2900), .clock(clock), .in1(R2899));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3101 (.out1(R3102), .clock(clock), .in1(R3101));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3348 (.out1(R3349), .clock(clock), .in1(R3348));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3540 (.out1(R3541), .clock(clock), .in1(R3540));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3728 (.out1(R3729), .clock(clock), .in1(R3728));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3945 (.out1(R3946), .clock(clock), .in1(_103));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3946 (.out1(R3947), .clock(clock), .in1(_164));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3947 (.out1(R3948), .clock(clock), .in1(_146));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3948 (.out1(R3949), .clock(clock), .in1(_139));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3949 (.out1(R3950), .clock(clock), .in1(_128));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3950 (.out1(R3951), .clock(clock), .in1(_121));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3951 (.out1(R3952), .clock(clock), .in1(_111));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3952 (.out1(R3953), .clock(clock), .in1(_104));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op104 (.out1(_96), .in1(R3349));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op155 (.out1(_147), .in1(R3948), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op173 (.out1(_165), .in1(R3947), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op156 (.out1(_148), .in1(R3949), .in2(_147));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op137 (.out1(_129), .in1(R3950), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op120 (.out1(_112), .in1(R3952), .in2(1 'd 1));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op138 (.out1(_130), .in1(R3951), .in2(_129));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op113 (.out1(_105), .in1(R3946), .in2(R3953));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op105 (.out1(_97), .in1(_96), .in2(2 'd 2));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op174 (.out1(_166), .in1(_165), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op157 (.out1(_149), .in1(_148), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op121 (.out1(_113), .in1(_112), .in2(63 'd 6148914691236517205));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op175 (.out1(_167), .in1(_149), .in2(_166));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op139 (.out1(_131), .in1(_130), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op122 (.out1(_114), .in1(_105), .in2(_113));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2694 (.out1(R2695), .clock(clock), .in1(R2694));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2900 (.out1(R2901), .clock(clock), .in1(R2900));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3102 (.out1(R3103), .clock(clock), .in1(R3102));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3349 (.out1(R3350), .clock(clock), .in1(R3349));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3541 (.out1(R3542), .clock(clock), .in1(R3541));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3729 (.out1(R3730), .clock(clock), .in1(R3729));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3953 (.out1(R3954), .clock(clock), .in1(_97));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3954 (.out1(R3955), .clock(clock), .in1(_167));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3955 (.out1(R3956), .clock(clock), .in1(_131));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3956 (.out1(R3957), .clock(clock), .in1(_114));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op140 (.out1(_132), .in1(R3956), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op123 (.out1(_115), .in1(R3957), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op176 (.out1(_168), .in1(R3955), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op141 (.out1(_133), .in1(_115), .in2(_132));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op106 (.out1(_98), .in1(c24_popcnt_2543_D), .in2(R3954));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op177 (.out1(_169), .in1(_133), .in2(_168));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op178 (.out1(_170), .in1(_169), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2695 (.out1(R2696), .clock(clock), .in1(R2695));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2901 (.out1(R2902), .clock(clock), .in1(R2901));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3103 (.out1(R3104), .clock(clock), .in1(R3103));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3350 (.out1(R3351), .clock(clock), .in1(R3350));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3542 (.out1(R3543), .clock(clock), .in1(R3542));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3730 (.out1(R3731), .clock(clock), .in1(R3730));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3957 (.out1(R3958), .clock(clock), .in1(_98));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3958 (.out1(R3959), .clock(clock), .in1(_170));
  SRAM op107 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_99),.ADR(R3958));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op179 (.out1(_171), .in1(R3959), .in2(57 'd 72340172838076673));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2696 (.out1(R2697), .clock(clock), .in1(R2696));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2902 (.out1(R2903), .clock(clock), .in1(R2902));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3104 (.out1(R3105), .clock(clock), .in1(R3104));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3351 (.out1(R3352), .clock(clock), .in1(R3351));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3543 (.out1(R3544), .clock(clock), .in1(R3543));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3731 (.out1(R3732), .clock(clock), .in1(R3731));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3959 (.out1(R3960), .clock(clock), .in1(_99));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3960 (.out1(R3961), .clock(clock), .in1(_171));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op180 (.out1(_172), .in1(R3961), .in2(6 'd 56));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op181 (.out1(_173), .in1(_172));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op182 (.out1(ck_idx_2544), .in1(R3960), .in2(_173));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2697 (.out1(R2698), .clock(clock), .in1(R2697));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2903 (.out1(R2904), .clock(clock), .in1(R2903));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3105 (.out1(R3106), .clock(clock), .in1(R3105));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3352 (.out1(R3353), .clock(clock), .in1(R3352));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3544 (.out1(R3545), .clock(clock), .in1(R3544));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3732 (.out1(R3733), .clock(clock), .in1(R3732));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3961 (.out1(R3962), .clock(clock), .in1(ck_idx_2544));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(4), .BITSIZE_out1(32), .PRECISION(32)) op183 (.out1(_174), .in1(R3962), .in2(4 'd 8));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op184 (.out1(_175), .in1(ip1_2522_D), .in2(6 'd 32));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2698 (.out1(R2699), .clock(clock), .in1(R2698));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2904 (.out1(R2905), .clock(clock), .in1(R2904));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3106 (.out1(R3107), .clock(clock), .in1(R3106));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3353 (.out1(R3354), .clock(clock), .in1(R3353));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3545 (.out1(R3546), .clock(clock), .in1(R3545));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3733 (.out1(R3734), .clock(clock), .in1(R3733));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3962 (.out1(R3963), .clock(clock), .in1(_174));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3963 (.out1(R3964), .clock(clock), .in1(_175));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op185 (.out1(_176), .in1(R3964));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(8), .BITSIZE_out1(32)) op186 (.out1(_177), .in1(_176), .in2(8 'd 255));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op187 (.out1(idx_sail_2545), .in1(R3963), .in2(_177));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(3), .BITSIZE_out1(32), .PRECISION(32)) op188 (.out1(idx_2546), .in1(idx_sail_2545), .in2(3 'd 6));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2699 (.out1(R2700), .clock(clock), .in1(R2699));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2905 (.out1(R2906), .clock(clock), .in1(R2905));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3107 (.out1(R3108), .clock(clock), .in1(R3107));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3354 (.out1(R3355), .clock(clock), .in1(R3354));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3546 (.out1(R3547), .clock(clock), .in1(R3546));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3734 (.out1(R3735), .clock(clock), .in1(R3734));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3964 (.out1(R3965), .clock(clock), .in1(idx_sail_2545));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3967 (.out1(R3968), .clock(clock), .in1(idx_2546));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op190 (.out1(_178), .in1(R3968));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op191 (.out1(_179), .in1(_178), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2700 (.out1(R2701), .clock(clock), .in1(R2700));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2906 (.out1(R2907), .clock(clock), .in1(R2906));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3108 (.out1(R3109), .clock(clock), .in1(R3108));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3355 (.out1(R3356), .clock(clock), .in1(R3355));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3547 (.out1(R3548), .clock(clock), .in1(R3547));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3735 (.out1(R3736), .clock(clock), .in1(R3735));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3965 (.out1(R3966), .clock(clock), .in1(R3965));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3968 (.out1(R3969), .clock(clock), .in1(R3968));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4145 (.out1(R4146), .clock(clock), .in1(_179));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op192 (.out1(_180), .in1(c32_bitmap_2548_D), .in2(R4146));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2701 (.out1(R2702), .clock(clock), .in1(R2701));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2907 (.out1(R2908), .clock(clock), .in1(R2907));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3109 (.out1(R3110), .clock(clock), .in1(R3109));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3356 (.out1(R3357), .clock(clock), .in1(R3356));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3548 (.out1(R3549), .clock(clock), .in1(R3548));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3736 (.out1(R3737), .clock(clock), .in1(R3736));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3966 (.out1(R3967), .clock(clock), .in1(R3966));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3969 (.out1(R3970), .clock(clock), .in1(R3969));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4146 (.out1(R4147), .clock(clock), .in1(_180));
  SRAM op193 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_181),.ADR(R4147));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op189 (.out1(off_2547), .in1(R3967), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op194 (.out1(_182), .in1(64 'd 9223372036854775808), .in2(off_2547));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2702 (.out1(R2703), .clock(clock), .in1(R2702));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2908 (.out1(R2909), .clock(clock), .in1(R2908));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3110 (.out1(R3111), .clock(clock), .in1(R3110));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3357 (.out1(R3358), .clock(clock), .in1(R3357));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3549 (.out1(R3550), .clock(clock), .in1(R3549));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3737 (.out1(R3738), .clock(clock), .in1(R3737));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3970 (.out1(R3971), .clock(clock), .in1(R3970));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4147 (.out1(R4148), .clock(clock), .in1(_181));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4148 (.out1(R4149), .clock(clock), .in1(off_2547));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4322 (.out1(R4323), .clock(clock), .in1(_182));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op195 (.out1(_183), .in1(R4148), .in2(R4323));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op196 (.out1(ifout196), .in1(_183), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op257 (.out1(_244), .in1(R3971));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op258 (.out1(_245), .in1(_244), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2703 (.out1(R2704), .clock(clock), .in1(R2703));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2909 (.out1(R2910), .clock(clock), .in1(R2909));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3111 (.out1(R3112), .clock(clock), .in1(R3111));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3358 (.out1(R3359), .clock(clock), .in1(R3358));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3550 (.out1(R3551), .clock(clock), .in1(R3550));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3738 (.out1(R3739), .clock(clock), .in1(R3738));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3971 (.out1(R3972), .clock(clock), .in1(R3971));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4149 (.out1(R4150), .clock(clock), .in1(R4149));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4323 (.out1(R4324), .clock(clock), .in1(ifout196));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4503 (.out1(R4504), .clock(clock), .in1(_245));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op251 (.out1(_238), .in1(R3972));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op241 (.out1(_228), .in1(R3972));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op235 (.out1(_222), .in1(R3972));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op223 (.out1(_210), .in1(R3972));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op217 (.out1(_204), .in1(R3972));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op207 (.out1(_194), .in1(R3972));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op252 (.out1(_239), .in1(_238), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op242 (.out1(_229), .in1(_228), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op236 (.out1(_223), .in1(_222), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op224 (.out1(_211), .in1(_210), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op218 (.out1(_205), .in1(_204), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op208 (.out1(_195), .in1(_194), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op259 (.out1(_246), .in1(c32_bitmap_2548_D), .in2(R4504));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2704 (.out1(R2705), .clock(clock), .in1(R2704));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2910 (.out1(R2911), .clock(clock), .in1(R2910));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3112 (.out1(R3113), .clock(clock), .in1(R3112));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3359 (.out1(R3360), .clock(clock), .in1(R3359));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3551 (.out1(R3552), .clock(clock), .in1(R3551));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3739 (.out1(R3740), .clock(clock), .in1(R3739));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3972 (.out1(R3973), .clock(clock), .in1(R3972));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4150 (.out1(R4151), .clock(clock), .in1(R4150));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4324 (.out1(R4325), .clock(clock), .in1(R4324));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4504 (.out1(R4505), .clock(clock), .in1(_239));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4505 (.out1(R4506), .clock(clock), .in1(_229));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4506 (.out1(R4507), .clock(clock), .in1(_223));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4507 (.out1(R4508), .clock(clock), .in1(_211));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4508 (.out1(R4509), .clock(clock), .in1(_205));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4509 (.out1(R4510), .clock(clock), .in1(_195));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4510 (.out1(R4511), .clock(clock), .in1(_246));
  SRAM op260 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_247),.ADR(R4511));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op201 (.out1(_188), .in1(R3973));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op202 (.out1(_189), .in1(_188), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op253 (.out1(_240), .in1(c32_bitmap_2548_D), .in2(R4505));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op243 (.out1(_230), .in1(c32_bitmap_2548_D), .in2(R4506));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op237 (.out1(_224), .in1(c32_bitmap_2548_D), .in2(R4507));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op225 (.out1(_212), .in1(c32_bitmap_2548_D), .in2(R4508));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op219 (.out1(_206), .in1(c32_bitmap_2548_D), .in2(R4509));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op209 (.out1(_196), .in1(c32_bitmap_2548_D), .in2(R4510));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2705 (.out1(R2706), .clock(clock), .in1(R2705));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2911 (.out1(R2912), .clock(clock), .in1(R2911));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3113 (.out1(R3114), .clock(clock), .in1(R3113));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3360 (.out1(R3361), .clock(clock), .in1(R3360));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3552 (.out1(R3553), .clock(clock), .in1(R3552));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3740 (.out1(R3741), .clock(clock), .in1(R3740));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3973 (.out1(R3974), .clock(clock), .in1(R3973));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4151 (.out1(R4152), .clock(clock), .in1(R4151));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4325 (.out1(R4326), .clock(clock), .in1(R4325));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4511 (.out1(R4512), .clock(clock), .in1(_247));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4512 (.out1(R4513), .clock(clock), .in1(_189));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4513 (.out1(R4514), .clock(clock), .in1(_240));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4514 (.out1(R4515), .clock(clock), .in1(_230));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4515 (.out1(R4516), .clock(clock), .in1(_224));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4516 (.out1(R4517), .clock(clock), .in1(_212));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4517 (.out1(R4518), .clock(clock), .in1(_206));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4518 (.out1(R4519), .clock(clock), .in1(_196));
  SRAM op254 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_241),.ADR(R4514));
  SRAM op244 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_231),.ADR(R4515));
  SRAM op238 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_225),.ADR(R4516));
  SRAM op226 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_213),.ADR(R4517));
  SRAM op220 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_207),.ADR(R4518));
  SRAM op210 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_197),.ADR(R4519));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op261 (.out1(_248), .in1(7 'd 64), .in2(R4152));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op203 (.out1(_190), .in1(c32_bitmap_2548_D), .in2(R4513));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op262 (.out1(_249), .in1(R4512), .in2(_248));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op255 (.out1(_242), .in1(7 'd 64), .in2(R4152));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op245 (.out1(_232), .in1(7 'd 64), .in2(R4152));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op227 (.out1(_214), .in1(7 'd 64), .in2(R4152));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2706 (.out1(R2707), .clock(clock), .in1(R2706));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2912 (.out1(R2913), .clock(clock), .in1(R2912));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3114 (.out1(R3115), .clock(clock), .in1(R3114));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3361 (.out1(R3362), .clock(clock), .in1(R3361));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3553 (.out1(R3554), .clock(clock), .in1(R3553));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3741 (.out1(R3742), .clock(clock), .in1(R3741));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3974 (.out1(R3975), .clock(clock), .in1(R3974));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4152 (.out1(R4153), .clock(clock), .in1(R4152));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4326 (.out1(R4327), .clock(clock), .in1(R4326));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4519 (.out1(R4520), .clock(clock), .in1(_241));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4520 (.out1(R4521), .clock(clock), .in1(_231));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4521 (.out1(R4522), .clock(clock), .in1(_225));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4522 (.out1(R4523), .clock(clock), .in1(_213));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4523 (.out1(R4524), .clock(clock), .in1(_207));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4524 (.out1(R4525), .clock(clock), .in1(_197));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4525 (.out1(R4526), .clock(clock), .in1(_190));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4526 (.out1(R4527), .clock(clock), .in1(_249));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4527 (.out1(R4528), .clock(clock), .in1(_242));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4528 (.out1(R4529), .clock(clock), .in1(_232));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4529 (.out1(R4530), .clock(clock), .in1(_214));
  SRAM op204 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_191),.ADR(R4526));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op263 (.out1(_250), .in1(R4527), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op256 (.out1(_243), .in1(R4520), .in2(R4528));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op246 (.out1(_233), .in1(R4521), .in2(R4529));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op239 (.out1(_226), .in1(7 'd 64), .in2(R4153));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op228 (.out1(_215), .in1(R4523), .in2(R4530));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op221 (.out1(_208), .in1(7 'd 64), .in2(R4153));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op211 (.out1(_198), .in1(7 'd 64), .in2(R4153));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op264 (.out1(_251), .in1(_250), .in2(63 'd 6148914691236517205));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op265 (.out1(_252), .in1(_243), .in2(_251));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op247 (.out1(_234), .in1(_233), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op240 (.out1(_227), .in1(R4522), .in2(_226));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op229 (.out1(_216), .in1(_215), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op222 (.out1(_209), .in1(R4524), .in2(_208));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op212 (.out1(_199), .in1(R4525), .in2(_198));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op205 (.out1(_192), .in1(7 'd 64), .in2(R4153));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2707 (.out1(R2708), .clock(clock), .in1(R2707));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2913 (.out1(R2914), .clock(clock), .in1(R2913));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3115 (.out1(R3116), .clock(clock), .in1(R3115));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3362 (.out1(R3363), .clock(clock), .in1(R3362));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3554 (.out1(R3555), .clock(clock), .in1(R3554));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3742 (.out1(R3743), .clock(clock), .in1(R3742));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3975 (.out1(R3976), .clock(clock), .in1(R3975));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4153 (.out1(R4154), .clock(clock), .in1(R4153));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4327 (.out1(R4328), .clock(clock), .in1(R4327));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4530 (.out1(R4531), .clock(clock), .in1(_191));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4531 (.out1(R4532), .clock(clock), .in1(_252));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4532 (.out1(R4533), .clock(clock), .in1(_234));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4533 (.out1(R4534), .clock(clock), .in1(_227));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4534 (.out1(R4535), .clock(clock), .in1(_216));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4535 (.out1(R4536), .clock(clock), .in1(_209));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4536 (.out1(R4537), .clock(clock), .in1(_199));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4537 (.out1(R4538), .clock(clock), .in1(_192));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op197 (.out1(_184), .in1(R3976));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op248 (.out1(_235), .in1(R4533), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op266 (.out1(_253), .in1(R4532), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op249 (.out1(_236), .in1(R4534), .in2(_235));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op230 (.out1(_217), .in1(R4535), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op213 (.out1(_200), .in1(R4537), .in2(1 'd 1));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op231 (.out1(_218), .in1(R4536), .in2(_217));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op206 (.out1(_193), .in1(R4531), .in2(R4538));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op198 (.out1(_185), .in1(_184), .in2(2 'd 2));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op267 (.out1(_254), .in1(_253), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op250 (.out1(_237), .in1(_236), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op214 (.out1(_201), .in1(_200), .in2(63 'd 6148914691236517205));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op268 (.out1(_255), .in1(_237), .in2(_254));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op232 (.out1(_219), .in1(_218), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op215 (.out1(_202), .in1(_193), .in2(_201));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2708 (.out1(R2709), .clock(clock), .in1(R2708));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2914 (.out1(R2915), .clock(clock), .in1(R2914));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3116 (.out1(R3117), .clock(clock), .in1(R3116));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3363 (.out1(R3364), .clock(clock), .in1(R3363));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3555 (.out1(R3556), .clock(clock), .in1(R3555));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3743 (.out1(R3744), .clock(clock), .in1(R3743));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3976 (.out1(R3977), .clock(clock), .in1(R3976));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4154 (.out1(R4155), .clock(clock), .in1(R4154));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4328 (.out1(R4329), .clock(clock), .in1(R4328));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4538 (.out1(R4539), .clock(clock), .in1(_185));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4539 (.out1(R4540), .clock(clock), .in1(_255));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4540 (.out1(R4541), .clock(clock), .in1(_219));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4541 (.out1(R4542), .clock(clock), .in1(_202));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op233 (.out1(_220), .in1(R4541), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op216 (.out1(_203), .in1(R4542), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op269 (.out1(_256), .in1(R4540), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op234 (.out1(_221), .in1(_203), .in2(_220));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op199 (.out1(_186), .in1(c32_popcnt_2553_D), .in2(R4539));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op270 (.out1(_257), .in1(_221), .in2(_256));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op271 (.out1(_258), .in1(_257), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2709 (.out1(R2710), .clock(clock), .in1(R2709));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2915 (.out1(R2916), .clock(clock), .in1(R2915));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3117 (.out1(R3118), .clock(clock), .in1(R3117));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3364 (.out1(R3365), .clock(clock), .in1(R3364));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3556 (.out1(R3557), .clock(clock), .in1(R3556));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3744 (.out1(R3745), .clock(clock), .in1(R3744));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3977 (.out1(R3978), .clock(clock), .in1(R3977));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4155 (.out1(R4156), .clock(clock), .in1(R4155));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4329 (.out1(R4330), .clock(clock), .in1(R4329));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4542 (.out1(R4543), .clock(clock), .in1(_186));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4543 (.out1(R4544), .clock(clock), .in1(_258));
  SRAM op200 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_187),.ADR(R4543));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op272 (.out1(_259), .in1(R4544), .in2(57 'd 72340172838076673));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2710 (.out1(R2711), .clock(clock), .in1(R2710));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2916 (.out1(R2917), .clock(clock), .in1(R2916));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3118 (.out1(R3119), .clock(clock), .in1(R3118));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3365 (.out1(R3366), .clock(clock), .in1(R3365));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3557 (.out1(R3558), .clock(clock), .in1(R3557));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3745 (.out1(R3746), .clock(clock), .in1(R3745));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3978 (.out1(R3979), .clock(clock), .in1(R3978));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4156 (.out1(R4157), .clock(clock), .in1(R4156));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4330 (.out1(R4331), .clock(clock), .in1(R4330));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4544 (.out1(R4545), .clock(clock), .in1(_187));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4545 (.out1(R4546), .clock(clock), .in1(_259));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op273 (.out1(_260), .in1(R4546), .in2(6 'd 56));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op274 (.out1(_261), .in1(_260));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op275 (.out1(ck_idx_2554), .in1(R4545), .in2(_261));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2711 (.out1(R2712), .clock(clock), .in1(R2711));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2917 (.out1(R2918), .clock(clock), .in1(R2917));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3119 (.out1(R3120), .clock(clock), .in1(R3119));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3366 (.out1(R3367), .clock(clock), .in1(R3366));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3558 (.out1(R3559), .clock(clock), .in1(R3558));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3746 (.out1(R3747), .clock(clock), .in1(R3746));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3979 (.out1(R3980), .clock(clock), .in1(R3979));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4157 (.out1(R4158), .clock(clock), .in1(R4157));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4331 (.out1(R4332), .clock(clock), .in1(R4331));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4546 (.out1(R4547), .clock(clock), .in1(ck_idx_2554));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(4), .BITSIZE_out1(32), .PRECISION(32)) op276 (.out1(_262), .in1(R4547), .in2(4 'd 8));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(5), .BITSIZE_out1(64), .PRECISION(64)) op277 (.out1(_263), .in1(ip1_2522_D), .in2(5 'd 24));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2712 (.out1(R2713), .clock(clock), .in1(R2712));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2918 (.out1(R2919), .clock(clock), .in1(R2918));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3120 (.out1(R3121), .clock(clock), .in1(R3120));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3367 (.out1(R3368), .clock(clock), .in1(R3367));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3559 (.out1(R3560), .clock(clock), .in1(R3559));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3747 (.out1(R3748), .clock(clock), .in1(R3747));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3980 (.out1(R3981), .clock(clock), .in1(R3980));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4158 (.out1(R4159), .clock(clock), .in1(R4158));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4332 (.out1(R4333), .clock(clock), .in1(R4332));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4547 (.out1(R4548), .clock(clock), .in1(_262));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4548 (.out1(R4549), .clock(clock), .in1(_263));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op278 (.out1(_264), .in1(R4549));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(8), .BITSIZE_out1(32)) op279 (.out1(_265), .in1(_264), .in2(8 'd 255));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op280 (.out1(idx_sail_2555), .in1(R4548), .in2(_265));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(3), .BITSIZE_out1(32), .PRECISION(32)) op281 (.out1(idx_2556), .in1(idx_sail_2555), .in2(3 'd 6));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2713 (.out1(R2714), .clock(clock), .in1(R2713));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2919 (.out1(R2920), .clock(clock), .in1(R2919));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3121 (.out1(R3122), .clock(clock), .in1(R3121));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3368 (.out1(R3369), .clock(clock), .in1(R3368));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3560 (.out1(R3561), .clock(clock), .in1(R3560));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3748 (.out1(R3749), .clock(clock), .in1(R3748));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3981 (.out1(R3982), .clock(clock), .in1(R3981));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4159 (.out1(R4160), .clock(clock), .in1(R4159));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4333 (.out1(R4334), .clock(clock), .in1(R4333));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4549 (.out1(R4550), .clock(clock), .in1(idx_sail_2555));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4552 (.out1(R4553), .clock(clock), .in1(idx_2556));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op283 (.out1(_266), .in1(R4553));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op284 (.out1(_267), .in1(_266), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2714 (.out1(R2715), .clock(clock), .in1(R2714));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2920 (.out1(R2921), .clock(clock), .in1(R2920));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3122 (.out1(R3123), .clock(clock), .in1(R3122));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3369 (.out1(R3370), .clock(clock), .in1(R3369));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3561 (.out1(R3562), .clock(clock), .in1(R3561));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3749 (.out1(R3750), .clock(clock), .in1(R3749));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3982 (.out1(R3983), .clock(clock), .in1(R3982));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4160 (.out1(R4161), .clock(clock), .in1(R4160));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4334 (.out1(R4335), .clock(clock), .in1(R4334));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4550 (.out1(R4551), .clock(clock), .in1(R4550));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4553 (.out1(R4554), .clock(clock), .in1(R4553));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4716 (.out1(R4717), .clock(clock), .in1(_267));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op285 (.out1(_268), .in1(c40_bitmap_2558_D), .in2(R4717));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2715 (.out1(R2716), .clock(clock), .in1(R2715));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2921 (.out1(R2922), .clock(clock), .in1(R2921));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3123 (.out1(R3124), .clock(clock), .in1(R3123));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3370 (.out1(R3371), .clock(clock), .in1(R3370));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3562 (.out1(R3563), .clock(clock), .in1(R3562));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3750 (.out1(R3751), .clock(clock), .in1(R3750));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3983 (.out1(R3984), .clock(clock), .in1(R3983));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4161 (.out1(R4162), .clock(clock), .in1(R4161));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4335 (.out1(R4336), .clock(clock), .in1(R4335));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4551 (.out1(R4552), .clock(clock), .in1(R4551));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4554 (.out1(R4555), .clock(clock), .in1(R4554));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4717 (.out1(R4718), .clock(clock), .in1(_268));
  SRAM op286 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_269),.ADR(R4718));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op282 (.out1(off_2557), .in1(R4552), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op287 (.out1(_270), .in1(64 'd 9223372036854775808), .in2(off_2557));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2716 (.out1(R2717), .clock(clock), .in1(R2716));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2922 (.out1(R2923), .clock(clock), .in1(R2922));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3124 (.out1(R3125), .clock(clock), .in1(R3124));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3371 (.out1(R3372), .clock(clock), .in1(R3371));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3563 (.out1(R3564), .clock(clock), .in1(R3563));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3751 (.out1(R3752), .clock(clock), .in1(R3751));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3984 (.out1(R3985), .clock(clock), .in1(R3984));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4162 (.out1(R4163), .clock(clock), .in1(R4162));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4336 (.out1(R4337), .clock(clock), .in1(R4336));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4555 (.out1(R4556), .clock(clock), .in1(R4555));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4718 (.out1(R4719), .clock(clock), .in1(_269));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4719 (.out1(R4720), .clock(clock), .in1(off_2557));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4879 (.out1(R4880), .clock(clock), .in1(_270));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op288 (.out1(_271), .in1(R4719), .in2(R4880));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op289 (.out1(ifout289), .in1(_271), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op350 (.out1(_332), .in1(R4556));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op351 (.out1(_333), .in1(_332), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2717 (.out1(R2718), .clock(clock), .in1(R2717));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2923 (.out1(R2924), .clock(clock), .in1(R2923));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3125 (.out1(R3126), .clock(clock), .in1(R3125));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3372 (.out1(R3373), .clock(clock), .in1(R3372));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3564 (.out1(R3565), .clock(clock), .in1(R3564));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3752 (.out1(R3753), .clock(clock), .in1(R3752));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3985 (.out1(R3986), .clock(clock), .in1(R3985));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4163 (.out1(R4164), .clock(clock), .in1(R4163));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4337 (.out1(R4338), .clock(clock), .in1(R4337));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4556 (.out1(R4557), .clock(clock), .in1(R4556));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4720 (.out1(R4721), .clock(clock), .in1(R4720));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4880 (.out1(R4881), .clock(clock), .in1(ifout289));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5046 (.out1(R5047), .clock(clock), .in1(_333));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op344 (.out1(_326), .in1(R4557));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op334 (.out1(_316), .in1(R4557));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op328 (.out1(_310), .in1(R4557));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op316 (.out1(_298), .in1(R4557));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op310 (.out1(_292), .in1(R4557));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op300 (.out1(_282), .in1(R4557));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op345 (.out1(_327), .in1(_326), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op335 (.out1(_317), .in1(_316), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op329 (.out1(_311), .in1(_310), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op317 (.out1(_299), .in1(_298), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op311 (.out1(_293), .in1(_292), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op301 (.out1(_283), .in1(_282), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op352 (.out1(_334), .in1(c40_bitmap_2558_D), .in2(R5047));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2718 (.out1(R2719), .clock(clock), .in1(R2718));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2924 (.out1(R2925), .clock(clock), .in1(R2924));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3126 (.out1(R3127), .clock(clock), .in1(R3126));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3373 (.out1(R3374), .clock(clock), .in1(R3373));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3565 (.out1(R3566), .clock(clock), .in1(R3565));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3753 (.out1(R3754), .clock(clock), .in1(R3753));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3986 (.out1(R3987), .clock(clock), .in1(R3986));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4164 (.out1(R4165), .clock(clock), .in1(R4164));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4338 (.out1(R4339), .clock(clock), .in1(R4338));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4557 (.out1(R4558), .clock(clock), .in1(R4557));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4721 (.out1(R4722), .clock(clock), .in1(R4721));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4881 (.out1(R4882), .clock(clock), .in1(R4881));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5047 (.out1(R5048), .clock(clock), .in1(_327));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5048 (.out1(R5049), .clock(clock), .in1(_317));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5049 (.out1(R5050), .clock(clock), .in1(_311));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5050 (.out1(R5051), .clock(clock), .in1(_299));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5051 (.out1(R5052), .clock(clock), .in1(_293));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5052 (.out1(R5053), .clock(clock), .in1(_283));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5053 (.out1(R5054), .clock(clock), .in1(_334));
  SRAM op353 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_335),.ADR(R5054));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op294 (.out1(_276), .in1(R4558));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op295 (.out1(_277), .in1(_276), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op346 (.out1(_328), .in1(c40_bitmap_2558_D), .in2(R5048));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op336 (.out1(_318), .in1(c40_bitmap_2558_D), .in2(R5049));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op330 (.out1(_312), .in1(c40_bitmap_2558_D), .in2(R5050));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op318 (.out1(_300), .in1(c40_bitmap_2558_D), .in2(R5051));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op312 (.out1(_294), .in1(c40_bitmap_2558_D), .in2(R5052));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op302 (.out1(_284), .in1(c40_bitmap_2558_D), .in2(R5053));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2719 (.out1(R2720), .clock(clock), .in1(R2719));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2925 (.out1(R2926), .clock(clock), .in1(R2925));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3127 (.out1(R3128), .clock(clock), .in1(R3127));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3374 (.out1(R3375), .clock(clock), .in1(R3374));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3566 (.out1(R3567), .clock(clock), .in1(R3566));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3754 (.out1(R3755), .clock(clock), .in1(R3754));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3987 (.out1(R3988), .clock(clock), .in1(R3987));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4165 (.out1(R4166), .clock(clock), .in1(R4165));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4339 (.out1(R4340), .clock(clock), .in1(R4339));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4558 (.out1(R4559), .clock(clock), .in1(R4558));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4722 (.out1(R4723), .clock(clock), .in1(R4722));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4882 (.out1(R4883), .clock(clock), .in1(R4882));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5054 (.out1(R5055), .clock(clock), .in1(_335));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5055 (.out1(R5056), .clock(clock), .in1(_277));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5056 (.out1(R5057), .clock(clock), .in1(_328));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5057 (.out1(R5058), .clock(clock), .in1(_318));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5058 (.out1(R5059), .clock(clock), .in1(_312));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5059 (.out1(R5060), .clock(clock), .in1(_300));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5060 (.out1(R5061), .clock(clock), .in1(_294));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5061 (.out1(R5062), .clock(clock), .in1(_284));
  SRAM op347 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_329),.ADR(R5057));
  SRAM op337 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_319),.ADR(R5058));
  SRAM op331 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_313),.ADR(R5059));
  SRAM op319 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_301),.ADR(R5060));
  SRAM op313 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_295),.ADR(R5061));
  SRAM op303 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_285),.ADR(R5062));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op354 (.out1(_336), .in1(7 'd 64), .in2(R4723));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op296 (.out1(_278), .in1(c40_bitmap_2558_D), .in2(R5056));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op355 (.out1(_337), .in1(R5055), .in2(_336));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op348 (.out1(_330), .in1(7 'd 64), .in2(R4723));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op338 (.out1(_320), .in1(7 'd 64), .in2(R4723));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op320 (.out1(_302), .in1(7 'd 64), .in2(R4723));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2720 (.out1(R2721), .clock(clock), .in1(R2720));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2926 (.out1(R2927), .clock(clock), .in1(R2926));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3128 (.out1(R3129), .clock(clock), .in1(R3128));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3375 (.out1(R3376), .clock(clock), .in1(R3375));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3567 (.out1(R3568), .clock(clock), .in1(R3567));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3755 (.out1(R3756), .clock(clock), .in1(R3755));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3988 (.out1(R3989), .clock(clock), .in1(R3988));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4166 (.out1(R4167), .clock(clock), .in1(R4166));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4340 (.out1(R4341), .clock(clock), .in1(R4340));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4559 (.out1(R4560), .clock(clock), .in1(R4559));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4723 (.out1(R4724), .clock(clock), .in1(R4723));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4883 (.out1(R4884), .clock(clock), .in1(R4883));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5062 (.out1(R5063), .clock(clock), .in1(_329));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5063 (.out1(R5064), .clock(clock), .in1(_319));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5064 (.out1(R5065), .clock(clock), .in1(_313));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5065 (.out1(R5066), .clock(clock), .in1(_301));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5066 (.out1(R5067), .clock(clock), .in1(_295));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5067 (.out1(R5068), .clock(clock), .in1(_285));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5068 (.out1(R5069), .clock(clock), .in1(_278));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5069 (.out1(R5070), .clock(clock), .in1(_337));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5070 (.out1(R5071), .clock(clock), .in1(_330));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5071 (.out1(R5072), .clock(clock), .in1(_320));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5072 (.out1(R5073), .clock(clock), .in1(_302));
  SRAM op297 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_279),.ADR(R5069));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op356 (.out1(_338), .in1(R5070), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op349 (.out1(_331), .in1(R5063), .in2(R5071));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op339 (.out1(_321), .in1(R5064), .in2(R5072));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op332 (.out1(_314), .in1(7 'd 64), .in2(R4724));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op321 (.out1(_303), .in1(R5066), .in2(R5073));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op314 (.out1(_296), .in1(7 'd 64), .in2(R4724));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op304 (.out1(_286), .in1(7 'd 64), .in2(R4724));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op357 (.out1(_339), .in1(_338), .in2(63 'd 6148914691236517205));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op358 (.out1(_340), .in1(_331), .in2(_339));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op340 (.out1(_322), .in1(_321), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op333 (.out1(_315), .in1(R5065), .in2(_314));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op322 (.out1(_304), .in1(_303), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op315 (.out1(_297), .in1(R5067), .in2(_296));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op305 (.out1(_287), .in1(R5068), .in2(_286));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op298 (.out1(_280), .in1(7 'd 64), .in2(R4724));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2721 (.out1(R2722), .clock(clock), .in1(R2721));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2927 (.out1(R2928), .clock(clock), .in1(R2927));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3129 (.out1(R3130), .clock(clock), .in1(R3129));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3376 (.out1(R3377), .clock(clock), .in1(R3376));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3568 (.out1(R3569), .clock(clock), .in1(R3568));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3756 (.out1(R3757), .clock(clock), .in1(R3756));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3989 (.out1(R3990), .clock(clock), .in1(R3989));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4167 (.out1(R4168), .clock(clock), .in1(R4167));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4341 (.out1(R4342), .clock(clock), .in1(R4341));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4560 (.out1(R4561), .clock(clock), .in1(R4560));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4724 (.out1(R4725), .clock(clock), .in1(R4724));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4884 (.out1(R4885), .clock(clock), .in1(R4884));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5073 (.out1(R5074), .clock(clock), .in1(_279));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5074 (.out1(R5075), .clock(clock), .in1(_340));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5075 (.out1(R5076), .clock(clock), .in1(_322));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5076 (.out1(R5077), .clock(clock), .in1(_315));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5077 (.out1(R5078), .clock(clock), .in1(_304));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5078 (.out1(R5079), .clock(clock), .in1(_297));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5079 (.out1(R5080), .clock(clock), .in1(_287));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5080 (.out1(R5081), .clock(clock), .in1(_280));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op290 (.out1(_272), .in1(R4561));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op341 (.out1(_323), .in1(R5076), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op359 (.out1(_341), .in1(R5075), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op342 (.out1(_324), .in1(R5077), .in2(_323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op323 (.out1(_305), .in1(R5078), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op306 (.out1(_288), .in1(R5080), .in2(1 'd 1));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op324 (.out1(_306), .in1(R5079), .in2(_305));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op299 (.out1(_281), .in1(R5074), .in2(R5081));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op291 (.out1(_273), .in1(_272), .in2(2 'd 2));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op360 (.out1(_342), .in1(_341), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op343 (.out1(_325), .in1(_324), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op307 (.out1(_289), .in1(_288), .in2(63 'd 6148914691236517205));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op361 (.out1(_343), .in1(_325), .in2(_342));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op325 (.out1(_307), .in1(_306), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op308 (.out1(_290), .in1(_281), .in2(_289));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2722 (.out1(R2723), .clock(clock), .in1(R2722));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2928 (.out1(R2929), .clock(clock), .in1(R2928));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3130 (.out1(R3131), .clock(clock), .in1(R3130));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3377 (.out1(R3378), .clock(clock), .in1(R3377));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3569 (.out1(R3570), .clock(clock), .in1(R3569));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3757 (.out1(R3758), .clock(clock), .in1(R3757));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3990 (.out1(R3991), .clock(clock), .in1(R3990));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4168 (.out1(R4169), .clock(clock), .in1(R4168));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4342 (.out1(R4343), .clock(clock), .in1(R4342));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4561 (.out1(R4562), .clock(clock), .in1(R4561));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4725 (.out1(R4726), .clock(clock), .in1(R4725));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4885 (.out1(R4886), .clock(clock), .in1(R4885));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5081 (.out1(R5082), .clock(clock), .in1(_273));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5082 (.out1(R5083), .clock(clock), .in1(_343));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5083 (.out1(R5084), .clock(clock), .in1(_307));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5084 (.out1(R5085), .clock(clock), .in1(_290));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op326 (.out1(_308), .in1(R5084), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op309 (.out1(_291), .in1(R5085), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op362 (.out1(_344), .in1(R5083), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op327 (.out1(_309), .in1(_291), .in2(_308));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op292 (.out1(_274), .in1(c40_popcnt_2563_D), .in2(R5082));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op363 (.out1(_345), .in1(_309), .in2(_344));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op364 (.out1(_346), .in1(_345), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2723 (.out1(R2724), .clock(clock), .in1(R2723));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2929 (.out1(R2930), .clock(clock), .in1(R2929));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3131 (.out1(R3132), .clock(clock), .in1(R3131));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3378 (.out1(R3379), .clock(clock), .in1(R3378));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3570 (.out1(R3571), .clock(clock), .in1(R3570));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3758 (.out1(R3759), .clock(clock), .in1(R3758));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3991 (.out1(R3992), .clock(clock), .in1(R3991));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4169 (.out1(R4170), .clock(clock), .in1(R4169));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4343 (.out1(R4344), .clock(clock), .in1(R4343));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4562 (.out1(R4563), .clock(clock), .in1(R4562));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4726 (.out1(R4727), .clock(clock), .in1(R4726));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4886 (.out1(R4887), .clock(clock), .in1(R4886));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5085 (.out1(R5086), .clock(clock), .in1(_274));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5086 (.out1(R5087), .clock(clock), .in1(_346));
  SRAM op293 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_275),.ADR(R5086));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op365 (.out1(_347), .in1(R5087), .in2(57 'd 72340172838076673));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2724 (.out1(R2725), .clock(clock), .in1(R2724));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2930 (.out1(R2931), .clock(clock), .in1(R2930));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3132 (.out1(R3133), .clock(clock), .in1(R3132));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3379 (.out1(R3380), .clock(clock), .in1(R3379));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3571 (.out1(R3572), .clock(clock), .in1(R3571));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3759 (.out1(R3760), .clock(clock), .in1(R3759));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3992 (.out1(R3993), .clock(clock), .in1(R3992));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4170 (.out1(R4171), .clock(clock), .in1(R4170));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4344 (.out1(R4345), .clock(clock), .in1(R4344));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4563 (.out1(R4564), .clock(clock), .in1(R4563));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4727 (.out1(R4728), .clock(clock), .in1(R4727));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4887 (.out1(R4888), .clock(clock), .in1(R4887));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5087 (.out1(R5088), .clock(clock), .in1(_275));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5088 (.out1(R5089), .clock(clock), .in1(_347));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op366 (.out1(_348), .in1(R5089), .in2(6 'd 56));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op367 (.out1(_349), .in1(_348));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op368 (.out1(ck_idx_2564), .in1(R5088), .in2(_349));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2725 (.out1(R2726), .clock(clock), .in1(R2725));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2931 (.out1(R2932), .clock(clock), .in1(R2931));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3133 (.out1(R3134), .clock(clock), .in1(R3133));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3380 (.out1(R3381), .clock(clock), .in1(R3380));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3572 (.out1(R3573), .clock(clock), .in1(R3572));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3760 (.out1(R3761), .clock(clock), .in1(R3760));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3993 (.out1(R3994), .clock(clock), .in1(R3993));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4171 (.out1(R4172), .clock(clock), .in1(R4171));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4345 (.out1(R4346), .clock(clock), .in1(R4345));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4564 (.out1(R4565), .clock(clock), .in1(R4564));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4728 (.out1(R4729), .clock(clock), .in1(R4728));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4888 (.out1(R4889), .clock(clock), .in1(R4888));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5089 (.out1(R5090), .clock(clock), .in1(ck_idx_2564));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(4), .BITSIZE_out1(32), .PRECISION(32)) op369 (.out1(_350), .in1(R5090), .in2(4 'd 8));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(5), .BITSIZE_out1(64), .PRECISION(64)) op370 (.out1(_351), .in1(ip1_2522_D), .in2(5 'd 16));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2726 (.out1(R2727), .clock(clock), .in1(R2726));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2932 (.out1(R2933), .clock(clock), .in1(R2932));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3134 (.out1(R3135), .clock(clock), .in1(R3134));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3381 (.out1(R3382), .clock(clock), .in1(R3381));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3573 (.out1(R3574), .clock(clock), .in1(R3573));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3761 (.out1(R3762), .clock(clock), .in1(R3761));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3994 (.out1(R3995), .clock(clock), .in1(R3994));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4172 (.out1(R4173), .clock(clock), .in1(R4172));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4346 (.out1(R4347), .clock(clock), .in1(R4346));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4565 (.out1(R4566), .clock(clock), .in1(R4565));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4729 (.out1(R4730), .clock(clock), .in1(R4729));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4889 (.out1(R4890), .clock(clock), .in1(R4889));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5090 (.out1(R5091), .clock(clock), .in1(_350));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5091 (.out1(R5092), .clock(clock), .in1(_351));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op371 (.out1(_352), .in1(R5092));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(8), .BITSIZE_out1(32)) op372 (.out1(_353), .in1(_352), .in2(8 'd 255));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op373 (.out1(idx_sail_2565), .in1(R5091), .in2(_353));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(3), .BITSIZE_out1(32), .PRECISION(32)) op374 (.out1(idx_2566), .in1(idx_sail_2565), .in2(3 'd 6));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2727 (.out1(R2728), .clock(clock), .in1(R2727));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2933 (.out1(R2934), .clock(clock), .in1(R2933));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3135 (.out1(R3136), .clock(clock), .in1(R3135));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3382 (.out1(R3383), .clock(clock), .in1(R3382));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3574 (.out1(R3575), .clock(clock), .in1(R3574));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3762 (.out1(R3763), .clock(clock), .in1(R3762));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3995 (.out1(R3996), .clock(clock), .in1(R3995));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4173 (.out1(R4174), .clock(clock), .in1(R4173));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4347 (.out1(R4348), .clock(clock), .in1(R4347));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4566 (.out1(R4567), .clock(clock), .in1(R4566));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4730 (.out1(R4731), .clock(clock), .in1(R4730));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4890 (.out1(R4891), .clock(clock), .in1(R4890));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5092 (.out1(R5093), .clock(clock), .in1(idx_sail_2565));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5095 (.out1(R5096), .clock(clock), .in1(idx_2566));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op376 (.out1(_354), .in1(R5096));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op377 (.out1(_355), .in1(_354), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2728 (.out1(R2729), .clock(clock), .in1(R2728));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2934 (.out1(R2935), .clock(clock), .in1(R2934));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3136 (.out1(R3137), .clock(clock), .in1(R3136));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3383 (.out1(R3384), .clock(clock), .in1(R3383));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3575 (.out1(R3576), .clock(clock), .in1(R3575));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3763 (.out1(R3764), .clock(clock), .in1(R3763));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3996 (.out1(R3997), .clock(clock), .in1(R3996));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4174 (.out1(R4175), .clock(clock), .in1(R4174));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4348 (.out1(R4349), .clock(clock), .in1(R4348));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4567 (.out1(R4568), .clock(clock), .in1(R4567));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4731 (.out1(R4732), .clock(clock), .in1(R4731));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4891 (.out1(R4892), .clock(clock), .in1(R4891));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5093 (.out1(R5094), .clock(clock), .in1(R5093));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5096 (.out1(R5097), .clock(clock), .in1(R5096));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5245 (.out1(R5246), .clock(clock), .in1(_355));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op378 (.out1(_356), .in1(c48_bitmap_2568_D), .in2(R5246));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2729 (.out1(R2730), .clock(clock), .in1(R2729));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2935 (.out1(R2936), .clock(clock), .in1(R2935));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3137 (.out1(R3138), .clock(clock), .in1(R3137));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3384 (.out1(R3385), .clock(clock), .in1(R3384));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3576 (.out1(R3577), .clock(clock), .in1(R3576));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3764 (.out1(R3765), .clock(clock), .in1(R3764));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3997 (.out1(R3998), .clock(clock), .in1(R3997));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4175 (.out1(R4176), .clock(clock), .in1(R4175));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4349 (.out1(R4350), .clock(clock), .in1(R4349));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4568 (.out1(R4569), .clock(clock), .in1(R4568));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4732 (.out1(R4733), .clock(clock), .in1(R4732));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4892 (.out1(R4893), .clock(clock), .in1(R4892));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5094 (.out1(R5095), .clock(clock), .in1(R5094));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5097 (.out1(R5098), .clock(clock), .in1(R5097));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5246 (.out1(R5247), .clock(clock), .in1(_356));
  SRAM op379 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_357),.ADR(R5247));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op375 (.out1(off_2567), .in1(R5095), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op380 (.out1(_358), .in1(64 'd 9223372036854775808), .in2(off_2567));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2730 (.out1(R2731), .clock(clock), .in1(R2730));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2936 (.out1(R2937), .clock(clock), .in1(R2936));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3138 (.out1(R3139), .clock(clock), .in1(R3138));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3385 (.out1(R3386), .clock(clock), .in1(R3385));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3577 (.out1(R3578), .clock(clock), .in1(R3577));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3765 (.out1(R3766), .clock(clock), .in1(R3765));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3998 (.out1(R3999), .clock(clock), .in1(R3998));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4176 (.out1(R4177), .clock(clock), .in1(R4176));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4350 (.out1(R4351), .clock(clock), .in1(R4350));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4569 (.out1(R4570), .clock(clock), .in1(R4569));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4733 (.out1(R4734), .clock(clock), .in1(R4733));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4893 (.out1(R4894), .clock(clock), .in1(R4893));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5098 (.out1(R5099), .clock(clock), .in1(R5098));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5247 (.out1(R5248), .clock(clock), .in1(_357));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5248 (.out1(R5249), .clock(clock), .in1(off_2567));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5394 (.out1(R5395), .clock(clock), .in1(_358));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op381 (.out1(_359), .in1(R5248), .in2(R5395));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op382 (.out1(ifout382), .in1(_359), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op443 (.out1(_420), .in1(R5099));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op444 (.out1(_421), .in1(_420), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2731 (.out1(R2732), .clock(clock), .in1(R2731));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2937 (.out1(R2938), .clock(clock), .in1(R2937));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3139 (.out1(R3140), .clock(clock), .in1(R3139));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3386 (.out1(R3387), .clock(clock), .in1(R3386));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3578 (.out1(R3579), .clock(clock), .in1(R3578));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3766 (.out1(R3767), .clock(clock), .in1(R3766));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3999 (.out1(R4000), .clock(clock), .in1(R3999));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4177 (.out1(R4178), .clock(clock), .in1(R4177));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4351 (.out1(R4352), .clock(clock), .in1(R4351));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4570 (.out1(R4571), .clock(clock), .in1(R4570));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4734 (.out1(R4735), .clock(clock), .in1(R4734));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4894 (.out1(R4895), .clock(clock), .in1(R4894));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5099 (.out1(R5100), .clock(clock), .in1(R5099));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5249 (.out1(R5250), .clock(clock), .in1(R5249));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5395 (.out1(R5396), .clock(clock), .in1(ifout382));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5547 (.out1(R5548), .clock(clock), .in1(_421));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op437 (.out1(_414), .in1(R5100));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op427 (.out1(_404), .in1(R5100));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op421 (.out1(_398), .in1(R5100));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op409 (.out1(_386), .in1(R5100));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op403 (.out1(_380), .in1(R5100));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op393 (.out1(_370), .in1(R5100));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op438 (.out1(_415), .in1(_414), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op428 (.out1(_405), .in1(_404), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op422 (.out1(_399), .in1(_398), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op410 (.out1(_387), .in1(_386), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op404 (.out1(_381), .in1(_380), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op394 (.out1(_371), .in1(_370), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op445 (.out1(_422), .in1(c48_bitmap_2568_D), .in2(R5548));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2732 (.out1(R2733), .clock(clock), .in1(R2732));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2938 (.out1(R2939), .clock(clock), .in1(R2938));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3140 (.out1(R3141), .clock(clock), .in1(R3140));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3387 (.out1(R3388), .clock(clock), .in1(R3387));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3579 (.out1(R3580), .clock(clock), .in1(R3579));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3767 (.out1(R3768), .clock(clock), .in1(R3767));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4000 (.out1(R4001), .clock(clock), .in1(R4000));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4178 (.out1(R4179), .clock(clock), .in1(R4178));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4352 (.out1(R4353), .clock(clock), .in1(R4352));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4571 (.out1(R4572), .clock(clock), .in1(R4571));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4735 (.out1(R4736), .clock(clock), .in1(R4735));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4895 (.out1(R4896), .clock(clock), .in1(R4895));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5100 (.out1(R5101), .clock(clock), .in1(R5100));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5250 (.out1(R5251), .clock(clock), .in1(R5250));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5396 (.out1(R5397), .clock(clock), .in1(R5396));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5548 (.out1(R5549), .clock(clock), .in1(_415));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5549 (.out1(R5550), .clock(clock), .in1(_405));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5550 (.out1(R5551), .clock(clock), .in1(_399));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5551 (.out1(R5552), .clock(clock), .in1(_387));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5552 (.out1(R5553), .clock(clock), .in1(_381));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5553 (.out1(R5554), .clock(clock), .in1(_371));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5554 (.out1(R5555), .clock(clock), .in1(_422));
  SRAM op446 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_423),.ADR(R5555));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op387 (.out1(_364), .in1(R5101));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op388 (.out1(_365), .in1(_364), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op439 (.out1(_416), .in1(c48_bitmap_2568_D), .in2(R5549));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op429 (.out1(_406), .in1(c48_bitmap_2568_D), .in2(R5550));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op423 (.out1(_400), .in1(c48_bitmap_2568_D), .in2(R5551));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op411 (.out1(_388), .in1(c48_bitmap_2568_D), .in2(R5552));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op405 (.out1(_382), .in1(c48_bitmap_2568_D), .in2(R5553));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op395 (.out1(_372), .in1(c48_bitmap_2568_D), .in2(R5554));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2733 (.out1(R2734), .clock(clock), .in1(R2733));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2939 (.out1(R2940), .clock(clock), .in1(R2939));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3141 (.out1(R3142), .clock(clock), .in1(R3141));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3388 (.out1(R3389), .clock(clock), .in1(R3388));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3580 (.out1(R3581), .clock(clock), .in1(R3580));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3768 (.out1(R3769), .clock(clock), .in1(R3768));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4001 (.out1(R4002), .clock(clock), .in1(R4001));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4179 (.out1(R4180), .clock(clock), .in1(R4179));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4353 (.out1(R4354), .clock(clock), .in1(R4353));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4572 (.out1(R4573), .clock(clock), .in1(R4572));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4736 (.out1(R4737), .clock(clock), .in1(R4736));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4896 (.out1(R4897), .clock(clock), .in1(R4896));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5101 (.out1(R5102), .clock(clock), .in1(R5101));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5251 (.out1(R5252), .clock(clock), .in1(R5251));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5397 (.out1(R5398), .clock(clock), .in1(R5397));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5555 (.out1(R5556), .clock(clock), .in1(_423));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5556 (.out1(R5557), .clock(clock), .in1(_365));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5557 (.out1(R5558), .clock(clock), .in1(_416));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5558 (.out1(R5559), .clock(clock), .in1(_406));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5559 (.out1(R5560), .clock(clock), .in1(_400));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5560 (.out1(R5561), .clock(clock), .in1(_388));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5561 (.out1(R5562), .clock(clock), .in1(_382));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5562 (.out1(R5563), .clock(clock), .in1(_372));
  SRAM op440 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_417),.ADR(R5558));
  SRAM op430 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_407),.ADR(R5559));
  SRAM op424 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_401),.ADR(R5560));
  SRAM op412 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_389),.ADR(R5561));
  SRAM op406 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_383),.ADR(R5562));
  SRAM op396 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_373),.ADR(R5563));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op447 (.out1(_424), .in1(7 'd 64), .in2(R5252));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op389 (.out1(_366), .in1(c48_bitmap_2568_D), .in2(R5557));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op448 (.out1(_425), .in1(R5556), .in2(_424));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op441 (.out1(_418), .in1(7 'd 64), .in2(R5252));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op431 (.out1(_408), .in1(7 'd 64), .in2(R5252));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op413 (.out1(_390), .in1(7 'd 64), .in2(R5252));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2734 (.out1(R2735), .clock(clock), .in1(R2734));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2940 (.out1(R2941), .clock(clock), .in1(R2940));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3142 (.out1(R3143), .clock(clock), .in1(R3142));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3389 (.out1(R3390), .clock(clock), .in1(R3389));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3581 (.out1(R3582), .clock(clock), .in1(R3581));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3769 (.out1(R3770), .clock(clock), .in1(R3769));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4002 (.out1(R4003), .clock(clock), .in1(R4002));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4180 (.out1(R4181), .clock(clock), .in1(R4180));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4354 (.out1(R4355), .clock(clock), .in1(R4354));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4573 (.out1(R4574), .clock(clock), .in1(R4573));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4737 (.out1(R4738), .clock(clock), .in1(R4737));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4897 (.out1(R4898), .clock(clock), .in1(R4897));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5102 (.out1(R5103), .clock(clock), .in1(R5102));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5252 (.out1(R5253), .clock(clock), .in1(R5252));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5398 (.out1(R5399), .clock(clock), .in1(R5398));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5563 (.out1(R5564), .clock(clock), .in1(_417));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5564 (.out1(R5565), .clock(clock), .in1(_407));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5565 (.out1(R5566), .clock(clock), .in1(_401));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5566 (.out1(R5567), .clock(clock), .in1(_389));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5567 (.out1(R5568), .clock(clock), .in1(_383));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5568 (.out1(R5569), .clock(clock), .in1(_373));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5569 (.out1(R5570), .clock(clock), .in1(_366));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5570 (.out1(R5571), .clock(clock), .in1(_425));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5571 (.out1(R5572), .clock(clock), .in1(_418));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5572 (.out1(R5573), .clock(clock), .in1(_408));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5573 (.out1(R5574), .clock(clock), .in1(_390));
  SRAM op390 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_367),.ADR(R5570));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op449 (.out1(_426), .in1(R5571), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op442 (.out1(_419), .in1(R5564), .in2(R5572));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op432 (.out1(_409), .in1(R5565), .in2(R5573));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op425 (.out1(_402), .in1(7 'd 64), .in2(R5253));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op414 (.out1(_391), .in1(R5567), .in2(R5574));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op407 (.out1(_384), .in1(7 'd 64), .in2(R5253));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op397 (.out1(_374), .in1(7 'd 64), .in2(R5253));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op450 (.out1(_427), .in1(_426), .in2(63 'd 6148914691236517205));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op451 (.out1(_428), .in1(_419), .in2(_427));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op433 (.out1(_410), .in1(_409), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op426 (.out1(_403), .in1(R5566), .in2(_402));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op415 (.out1(_392), .in1(_391), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op408 (.out1(_385), .in1(R5568), .in2(_384));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op398 (.out1(_375), .in1(R5569), .in2(_374));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op391 (.out1(_368), .in1(7 'd 64), .in2(R5253));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2735 (.out1(R2736), .clock(clock), .in1(R2735));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2941 (.out1(R2942), .clock(clock), .in1(R2941));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3143 (.out1(R3144), .clock(clock), .in1(R3143));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3390 (.out1(R3391), .clock(clock), .in1(R3390));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3582 (.out1(R3583), .clock(clock), .in1(R3582));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3770 (.out1(R3771), .clock(clock), .in1(R3770));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4003 (.out1(R4004), .clock(clock), .in1(R4003));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4181 (.out1(R4182), .clock(clock), .in1(R4181));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4355 (.out1(R4356), .clock(clock), .in1(R4355));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4574 (.out1(R4575), .clock(clock), .in1(R4574));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4738 (.out1(R4739), .clock(clock), .in1(R4738));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4898 (.out1(R4899), .clock(clock), .in1(R4898));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5103 (.out1(R5104), .clock(clock), .in1(R5103));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5253 (.out1(R5254), .clock(clock), .in1(R5253));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5399 (.out1(R5400), .clock(clock), .in1(R5399));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5574 (.out1(R5575), .clock(clock), .in1(_367));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5575 (.out1(R5576), .clock(clock), .in1(_428));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5576 (.out1(R5577), .clock(clock), .in1(_410));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5577 (.out1(R5578), .clock(clock), .in1(_403));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5578 (.out1(R5579), .clock(clock), .in1(_392));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5579 (.out1(R5580), .clock(clock), .in1(_385));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5580 (.out1(R5581), .clock(clock), .in1(_375));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5581 (.out1(R5582), .clock(clock), .in1(_368));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op383 (.out1(_360), .in1(R5104));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op434 (.out1(_411), .in1(R5577), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op452 (.out1(_429), .in1(R5576), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op435 (.out1(_412), .in1(R5578), .in2(_411));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op416 (.out1(_393), .in1(R5579), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op399 (.out1(_376), .in1(R5581), .in2(1 'd 1));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op417 (.out1(_394), .in1(R5580), .in2(_393));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op392 (.out1(_369), .in1(R5575), .in2(R5582));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op384 (.out1(_361), .in1(_360), .in2(2 'd 2));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op453 (.out1(_430), .in1(_429), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op436 (.out1(_413), .in1(_412), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op400 (.out1(_377), .in1(_376), .in2(63 'd 6148914691236517205));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op454 (.out1(_431), .in1(_413), .in2(_430));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op418 (.out1(_395), .in1(_394), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op401 (.out1(_378), .in1(_369), .in2(_377));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2736 (.out1(R2737), .clock(clock), .in1(R2736));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2942 (.out1(R2943), .clock(clock), .in1(R2942));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3144 (.out1(R3145), .clock(clock), .in1(R3144));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3391 (.out1(R3392), .clock(clock), .in1(R3391));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3583 (.out1(R3584), .clock(clock), .in1(R3583));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3771 (.out1(R3772), .clock(clock), .in1(R3771));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4004 (.out1(R4005), .clock(clock), .in1(R4004));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4182 (.out1(R4183), .clock(clock), .in1(R4182));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4356 (.out1(R4357), .clock(clock), .in1(R4356));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4575 (.out1(R4576), .clock(clock), .in1(R4575));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4739 (.out1(R4740), .clock(clock), .in1(R4739));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4899 (.out1(R4900), .clock(clock), .in1(R4899));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5104 (.out1(R5105), .clock(clock), .in1(R5104));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5254 (.out1(R5255), .clock(clock), .in1(R5254));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5400 (.out1(R5401), .clock(clock), .in1(R5400));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5582 (.out1(R5583), .clock(clock), .in1(_361));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5583 (.out1(R5584), .clock(clock), .in1(_431));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5584 (.out1(R5585), .clock(clock), .in1(_395));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5585 (.out1(R5586), .clock(clock), .in1(_378));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op419 (.out1(_396), .in1(R5585), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op402 (.out1(_379), .in1(R5586), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op455 (.out1(_432), .in1(R5584), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op420 (.out1(_397), .in1(_379), .in2(_396));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op385 (.out1(_362), .in1(c48_popcnt_2573_D), .in2(R5583));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op456 (.out1(_433), .in1(_397), .in2(_432));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op457 (.out1(_434), .in1(_433), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2737 (.out1(R2738), .clock(clock), .in1(R2737));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2943 (.out1(R2944), .clock(clock), .in1(R2943));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3145 (.out1(R3146), .clock(clock), .in1(R3145));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3392 (.out1(R3393), .clock(clock), .in1(R3392));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3584 (.out1(R3585), .clock(clock), .in1(R3584));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3772 (.out1(R3773), .clock(clock), .in1(R3772));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4005 (.out1(R4006), .clock(clock), .in1(R4005));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4183 (.out1(R4184), .clock(clock), .in1(R4183));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4357 (.out1(R4358), .clock(clock), .in1(R4357));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4576 (.out1(R4577), .clock(clock), .in1(R4576));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4740 (.out1(R4741), .clock(clock), .in1(R4740));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4900 (.out1(R4901), .clock(clock), .in1(R4900));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5105 (.out1(R5106), .clock(clock), .in1(R5105));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5255 (.out1(R5256), .clock(clock), .in1(R5255));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5401 (.out1(R5402), .clock(clock), .in1(R5401));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5586 (.out1(R5587), .clock(clock), .in1(_362));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5587 (.out1(R5588), .clock(clock), .in1(_434));
  SRAM op386 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_363),.ADR(R5587));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op458 (.out1(_435), .in1(R5588), .in2(57 'd 72340172838076673));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2738 (.out1(R2739), .clock(clock), .in1(R2738));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2944 (.out1(R2945), .clock(clock), .in1(R2944));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3146 (.out1(R3147), .clock(clock), .in1(R3146));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3393 (.out1(R3394), .clock(clock), .in1(R3393));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3585 (.out1(R3586), .clock(clock), .in1(R3585));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3773 (.out1(R3774), .clock(clock), .in1(R3773));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4006 (.out1(R4007), .clock(clock), .in1(R4006));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4184 (.out1(R4185), .clock(clock), .in1(R4184));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4358 (.out1(R4359), .clock(clock), .in1(R4358));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4577 (.out1(R4578), .clock(clock), .in1(R4577));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4741 (.out1(R4742), .clock(clock), .in1(R4741));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4901 (.out1(R4902), .clock(clock), .in1(R4901));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5106 (.out1(R5107), .clock(clock), .in1(R5106));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5256 (.out1(R5257), .clock(clock), .in1(R5256));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5402 (.out1(R5403), .clock(clock), .in1(R5402));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5588 (.out1(R5589), .clock(clock), .in1(_363));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5589 (.out1(R5590), .clock(clock), .in1(_435));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op459 (.out1(_436), .in1(R5590), .in2(6 'd 56));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op460 (.out1(_437), .in1(_436));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op461 (.out1(ck_idx_2574), .in1(R5589), .in2(_437));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2739 (.out1(R2740), .clock(clock), .in1(R2739));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2945 (.out1(R2946), .clock(clock), .in1(R2945));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3147 (.out1(R3148), .clock(clock), .in1(R3147));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3394 (.out1(R3395), .clock(clock), .in1(R3394));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3586 (.out1(R3587), .clock(clock), .in1(R3586));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3774 (.out1(R3775), .clock(clock), .in1(R3774));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4007 (.out1(R4008), .clock(clock), .in1(R4007));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4185 (.out1(R4186), .clock(clock), .in1(R4185));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4359 (.out1(R4360), .clock(clock), .in1(R4359));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4578 (.out1(R4579), .clock(clock), .in1(R4578));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4742 (.out1(R4743), .clock(clock), .in1(R4742));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4902 (.out1(R4903), .clock(clock), .in1(R4902));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5107 (.out1(R5108), .clock(clock), .in1(R5107));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5257 (.out1(R5258), .clock(clock), .in1(R5257));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5403 (.out1(R5404), .clock(clock), .in1(R5403));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5590 (.out1(R5591), .clock(clock), .in1(ck_idx_2574));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(4), .BITSIZE_out1(32), .PRECISION(32)) op462 (.out1(_438), .in1(R5591), .in2(4 'd 8));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(4), .BITSIZE_out1(64), .PRECISION(64)) op463 (.out1(_439), .in1(ip1_2522_D), .in2(4 'd 8));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2740 (.out1(R2741), .clock(clock), .in1(R2740));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2946 (.out1(R2947), .clock(clock), .in1(R2946));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3148 (.out1(R3149), .clock(clock), .in1(R3148));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3395 (.out1(R3396), .clock(clock), .in1(R3395));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3587 (.out1(R3588), .clock(clock), .in1(R3587));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3775 (.out1(R3776), .clock(clock), .in1(R3775));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4008 (.out1(R4009), .clock(clock), .in1(R4008));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4186 (.out1(R4187), .clock(clock), .in1(R4186));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4360 (.out1(R4361), .clock(clock), .in1(R4360));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4579 (.out1(R4580), .clock(clock), .in1(R4579));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4743 (.out1(R4744), .clock(clock), .in1(R4743));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4903 (.out1(R4904), .clock(clock), .in1(R4903));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5108 (.out1(R5109), .clock(clock), .in1(R5108));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5258 (.out1(R5259), .clock(clock), .in1(R5258));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5404 (.out1(R5405), .clock(clock), .in1(R5404));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5591 (.out1(R5592), .clock(clock), .in1(_438));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5592 (.out1(R5593), .clock(clock), .in1(_439));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op464 (.out1(_440), .in1(R5593));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(8), .BITSIZE_out1(32)) op465 (.out1(_441), .in1(_440), .in2(8 'd 255));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op466 (.out1(idx_sail_2575), .in1(R5592), .in2(_441));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(3), .BITSIZE_out1(32), .PRECISION(32)) op467 (.out1(idx_2576), .in1(idx_sail_2575), .in2(3 'd 6));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2741 (.out1(R2742), .clock(clock), .in1(R2741));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2947 (.out1(R2948), .clock(clock), .in1(R2947));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3149 (.out1(R3150), .clock(clock), .in1(R3149));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3396 (.out1(R3397), .clock(clock), .in1(R3396));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3588 (.out1(R3589), .clock(clock), .in1(R3588));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3776 (.out1(R3777), .clock(clock), .in1(R3776));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4009 (.out1(R4010), .clock(clock), .in1(R4009));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4187 (.out1(R4188), .clock(clock), .in1(R4187));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4361 (.out1(R4362), .clock(clock), .in1(R4361));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4580 (.out1(R4581), .clock(clock), .in1(R4580));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4744 (.out1(R4745), .clock(clock), .in1(R4744));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4904 (.out1(R4905), .clock(clock), .in1(R4904));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5109 (.out1(R5110), .clock(clock), .in1(R5109));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5259 (.out1(R5260), .clock(clock), .in1(R5259));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5405 (.out1(R5406), .clock(clock), .in1(R5405));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5593 (.out1(R5594), .clock(clock), .in1(idx_sail_2575));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5596 (.out1(R5597), .clock(clock), .in1(idx_2576));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op469 (.out1(_442), .in1(R5597));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op470 (.out1(_443), .in1(_442), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2742 (.out1(R2743), .clock(clock), .in1(R2742));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2948 (.out1(R2949), .clock(clock), .in1(R2948));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3150 (.out1(R3151), .clock(clock), .in1(R3150));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3397 (.out1(R3398), .clock(clock), .in1(R3397));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3589 (.out1(R3590), .clock(clock), .in1(R3589));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3777 (.out1(R3778), .clock(clock), .in1(R3777));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4010 (.out1(R4011), .clock(clock), .in1(R4010));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4188 (.out1(R4189), .clock(clock), .in1(R4188));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4362 (.out1(R4363), .clock(clock), .in1(R4362));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4581 (.out1(R4582), .clock(clock), .in1(R4581));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4745 (.out1(R4746), .clock(clock), .in1(R4745));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4905 (.out1(R4906), .clock(clock), .in1(R4905));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5110 (.out1(R5111), .clock(clock), .in1(R5110));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5260 (.out1(R5261), .clock(clock), .in1(R5260));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5406 (.out1(R5407), .clock(clock), .in1(R5406));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5594 (.out1(R5595), .clock(clock), .in1(R5594));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5597 (.out1(R5598), .clock(clock), .in1(R5597));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5732 (.out1(R5733), .clock(clock), .in1(_443));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op471 (.out1(_444), .in1(c56_bitmap_2578_D), .in2(R5733));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2743 (.out1(R2744), .clock(clock), .in1(R2743));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2949 (.out1(R2950), .clock(clock), .in1(R2949));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3151 (.out1(R3152), .clock(clock), .in1(R3151));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3398 (.out1(R3399), .clock(clock), .in1(R3398));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3590 (.out1(R3591), .clock(clock), .in1(R3590));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3778 (.out1(R3779), .clock(clock), .in1(R3778));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4011 (.out1(R4012), .clock(clock), .in1(R4011));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4189 (.out1(R4190), .clock(clock), .in1(R4189));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4363 (.out1(R4364), .clock(clock), .in1(R4363));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4582 (.out1(R4583), .clock(clock), .in1(R4582));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4746 (.out1(R4747), .clock(clock), .in1(R4746));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4906 (.out1(R4907), .clock(clock), .in1(R4906));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5111 (.out1(R5112), .clock(clock), .in1(R5111));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5261 (.out1(R5262), .clock(clock), .in1(R5261));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5407 (.out1(R5408), .clock(clock), .in1(R5407));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5595 (.out1(R5596), .clock(clock), .in1(R5595));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5598 (.out1(R5599), .clock(clock), .in1(R5598));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5733 (.out1(R5734), .clock(clock), .in1(_444));
  SRAM op472 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_445),.ADR(R5734));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op468 (.out1(off_2577), .in1(R5596), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op473 (.out1(_446), .in1(64 'd 9223372036854775808), .in2(off_2577));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2744 (.out1(R2745), .clock(clock), .in1(R2744));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2950 (.out1(R2951), .clock(clock), .in1(R2950));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3152 (.out1(R3153), .clock(clock), .in1(R3152));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3399 (.out1(R3400), .clock(clock), .in1(R3399));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3591 (.out1(R3592), .clock(clock), .in1(R3591));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3779 (.out1(R3780), .clock(clock), .in1(R3779));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4012 (.out1(R4013), .clock(clock), .in1(R4012));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4190 (.out1(R4191), .clock(clock), .in1(R4190));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4364 (.out1(R4365), .clock(clock), .in1(R4364));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4583 (.out1(R4584), .clock(clock), .in1(R4583));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4747 (.out1(R4748), .clock(clock), .in1(R4747));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4907 (.out1(R4908), .clock(clock), .in1(R4907));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5112 (.out1(R5113), .clock(clock), .in1(R5112));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5262 (.out1(R5263), .clock(clock), .in1(R5262));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5408 (.out1(R5409), .clock(clock), .in1(R5408));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5599 (.out1(R5600), .clock(clock), .in1(R5599));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5734 (.out1(R5735), .clock(clock), .in1(_445));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5735 (.out1(R5736), .clock(clock), .in1(off_2577));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5867 (.out1(R5868), .clock(clock), .in1(_446));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op474 (.out1(_447), .in1(R5735), .in2(R5868));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op475 (.out1(ifout475), .in1(_447), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op536 (.out1(_508), .in1(R5600));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op537 (.out1(_509), .in1(_508), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2745 (.out1(R2746), .clock(clock), .in1(R2745));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2951 (.out1(R2952), .clock(clock), .in1(R2951));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3153 (.out1(R3154), .clock(clock), .in1(R3153));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3400 (.out1(R3401), .clock(clock), .in1(R3400));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3592 (.out1(R3593), .clock(clock), .in1(R3592));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3780 (.out1(R3781), .clock(clock), .in1(R3780));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4013 (.out1(R4014), .clock(clock), .in1(R4013));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4191 (.out1(R4192), .clock(clock), .in1(R4191));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4365 (.out1(R4366), .clock(clock), .in1(R4365));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4584 (.out1(R4585), .clock(clock), .in1(R4584));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4748 (.out1(R4749), .clock(clock), .in1(R4748));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4908 (.out1(R4909), .clock(clock), .in1(R4908));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5113 (.out1(R5114), .clock(clock), .in1(R5113));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5263 (.out1(R5264), .clock(clock), .in1(R5263));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5409 (.out1(R5410), .clock(clock), .in1(R5409));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5600 (.out1(R5601), .clock(clock), .in1(R5600));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5736 (.out1(R5737), .clock(clock), .in1(R5736));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5868 (.out1(R5869), .clock(clock), .in1(ifout475));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6006 (.out1(R6007), .clock(clock), .in1(_509));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op530 (.out1(_502), .in1(R5601));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op520 (.out1(_492), .in1(R5601));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op514 (.out1(_486), .in1(R5601));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op502 (.out1(_474), .in1(R5601));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op496 (.out1(_468), .in1(R5601));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op486 (.out1(_458), .in1(R5601));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op531 (.out1(_503), .in1(_502), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op521 (.out1(_493), .in1(_492), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op515 (.out1(_487), .in1(_486), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op503 (.out1(_475), .in1(_474), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op497 (.out1(_469), .in1(_468), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op487 (.out1(_459), .in1(_458), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op538 (.out1(_510), .in1(c56_bitmap_2578_D), .in2(R6007));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2746 (.out1(R2747), .clock(clock), .in1(R2746));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2952 (.out1(R2953), .clock(clock), .in1(R2952));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3154 (.out1(R3155), .clock(clock), .in1(R3154));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3401 (.out1(R3402), .clock(clock), .in1(R3401));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3593 (.out1(R3594), .clock(clock), .in1(R3593));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3781 (.out1(R3782), .clock(clock), .in1(R3781));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4014 (.out1(R4015), .clock(clock), .in1(R4014));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4192 (.out1(R4193), .clock(clock), .in1(R4192));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4366 (.out1(R4367), .clock(clock), .in1(R4366));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4585 (.out1(R4586), .clock(clock), .in1(R4585));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4749 (.out1(R4750), .clock(clock), .in1(R4749));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4909 (.out1(R4910), .clock(clock), .in1(R4909));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5114 (.out1(R5115), .clock(clock), .in1(R5114));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5264 (.out1(R5265), .clock(clock), .in1(R5264));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5410 (.out1(R5411), .clock(clock), .in1(R5410));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5601 (.out1(R5602), .clock(clock), .in1(R5601));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5737 (.out1(R5738), .clock(clock), .in1(R5737));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5869 (.out1(R5870), .clock(clock), .in1(R5869));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6007 (.out1(R6008), .clock(clock), .in1(_503));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6008 (.out1(R6009), .clock(clock), .in1(_493));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6009 (.out1(R6010), .clock(clock), .in1(_487));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6010 (.out1(R6011), .clock(clock), .in1(_475));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6011 (.out1(R6012), .clock(clock), .in1(_469));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6012 (.out1(R6013), .clock(clock), .in1(_459));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6013 (.out1(R6014), .clock(clock), .in1(_510));
  SRAM op539 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_511),.ADR(R6014));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op480 (.out1(_452), .in1(R5602));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op481 (.out1(_453), .in1(_452), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op532 (.out1(_504), .in1(c56_bitmap_2578_D), .in2(R6008));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op522 (.out1(_494), .in1(c56_bitmap_2578_D), .in2(R6009));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op516 (.out1(_488), .in1(c56_bitmap_2578_D), .in2(R6010));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op504 (.out1(_476), .in1(c56_bitmap_2578_D), .in2(R6011));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op498 (.out1(_470), .in1(c56_bitmap_2578_D), .in2(R6012));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op488 (.out1(_460), .in1(c56_bitmap_2578_D), .in2(R6013));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2747 (.out1(R2748), .clock(clock), .in1(R2747));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2953 (.out1(R2954), .clock(clock), .in1(R2953));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3155 (.out1(R3156), .clock(clock), .in1(R3155));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3402 (.out1(R3403), .clock(clock), .in1(R3402));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3594 (.out1(R3595), .clock(clock), .in1(R3594));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3782 (.out1(R3783), .clock(clock), .in1(R3782));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4015 (.out1(R4016), .clock(clock), .in1(R4015));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4193 (.out1(R4194), .clock(clock), .in1(R4193));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4367 (.out1(R4368), .clock(clock), .in1(R4367));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4586 (.out1(R4587), .clock(clock), .in1(R4586));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4750 (.out1(R4751), .clock(clock), .in1(R4750));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4910 (.out1(R4911), .clock(clock), .in1(R4910));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5115 (.out1(R5116), .clock(clock), .in1(R5115));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5265 (.out1(R5266), .clock(clock), .in1(R5265));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5411 (.out1(R5412), .clock(clock), .in1(R5411));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5602 (.out1(R5603), .clock(clock), .in1(R5602));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5738 (.out1(R5739), .clock(clock), .in1(R5738));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5870 (.out1(R5871), .clock(clock), .in1(R5870));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6014 (.out1(R6015), .clock(clock), .in1(_511));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6015 (.out1(R6016), .clock(clock), .in1(_453));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6016 (.out1(R6017), .clock(clock), .in1(_504));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6017 (.out1(R6018), .clock(clock), .in1(_494));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6018 (.out1(R6019), .clock(clock), .in1(_488));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6019 (.out1(R6020), .clock(clock), .in1(_476));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6020 (.out1(R6021), .clock(clock), .in1(_470));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6021 (.out1(R6022), .clock(clock), .in1(_460));
  SRAM op533 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_505),.ADR(R6017));
  SRAM op523 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_495),.ADR(R6018));
  SRAM op517 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_489),.ADR(R6019));
  SRAM op505 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_477),.ADR(R6020));
  SRAM op499 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_471),.ADR(R6021));
  SRAM op489 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_461),.ADR(R6022));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op540 (.out1(_512), .in1(7 'd 64), .in2(R5739));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op482 (.out1(_454), .in1(c56_bitmap_2578_D), .in2(R6016));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op541 (.out1(_513), .in1(R6015), .in2(_512));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op534 (.out1(_506), .in1(7 'd 64), .in2(R5739));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op524 (.out1(_496), .in1(7 'd 64), .in2(R5739));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op506 (.out1(_478), .in1(7 'd 64), .in2(R5739));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2748 (.out1(R2749), .clock(clock), .in1(R2748));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2954 (.out1(R2955), .clock(clock), .in1(R2954));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3156 (.out1(R3157), .clock(clock), .in1(R3156));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3403 (.out1(R3404), .clock(clock), .in1(R3403));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3595 (.out1(R3596), .clock(clock), .in1(R3595));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3783 (.out1(R3784), .clock(clock), .in1(R3783));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4016 (.out1(R4017), .clock(clock), .in1(R4016));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4194 (.out1(R4195), .clock(clock), .in1(R4194));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4368 (.out1(R4369), .clock(clock), .in1(R4368));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4587 (.out1(R4588), .clock(clock), .in1(R4587));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4751 (.out1(R4752), .clock(clock), .in1(R4751));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4911 (.out1(R4912), .clock(clock), .in1(R4911));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5116 (.out1(R5117), .clock(clock), .in1(R5116));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5266 (.out1(R5267), .clock(clock), .in1(R5266));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5412 (.out1(R5413), .clock(clock), .in1(R5412));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5603 (.out1(R5604), .clock(clock), .in1(R5603));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5739 (.out1(R5740), .clock(clock), .in1(R5739));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5871 (.out1(R5872), .clock(clock), .in1(R5871));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6022 (.out1(R6023), .clock(clock), .in1(_505));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6023 (.out1(R6024), .clock(clock), .in1(_495));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6024 (.out1(R6025), .clock(clock), .in1(_489));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6025 (.out1(R6026), .clock(clock), .in1(_477));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6026 (.out1(R6027), .clock(clock), .in1(_471));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6027 (.out1(R6028), .clock(clock), .in1(_461));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6028 (.out1(R6029), .clock(clock), .in1(_454));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6029 (.out1(R6030), .clock(clock), .in1(_513));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6030 (.out1(R6031), .clock(clock), .in1(_506));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6031 (.out1(R6032), .clock(clock), .in1(_496));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6032 (.out1(R6033), .clock(clock), .in1(_478));
  SRAM op483 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_455),.ADR(R6029));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op542 (.out1(_514), .in1(R6030), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op535 (.out1(_507), .in1(R6023), .in2(R6031));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op525 (.out1(_497), .in1(R6024), .in2(R6032));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op518 (.out1(_490), .in1(7 'd 64), .in2(R5740));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op507 (.out1(_479), .in1(R6026), .in2(R6033));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op500 (.out1(_472), .in1(7 'd 64), .in2(R5740));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op490 (.out1(_462), .in1(7 'd 64), .in2(R5740));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op543 (.out1(_515), .in1(_514), .in2(63 'd 6148914691236517205));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op544 (.out1(_516), .in1(_507), .in2(_515));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op526 (.out1(_498), .in1(_497), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op519 (.out1(_491), .in1(R6025), .in2(_490));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op508 (.out1(_480), .in1(_479), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op501 (.out1(_473), .in1(R6027), .in2(_472));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op491 (.out1(_463), .in1(R6028), .in2(_462));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op484 (.out1(_456), .in1(7 'd 64), .in2(R5740));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2749 (.out1(R2750), .clock(clock), .in1(R2749));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2955 (.out1(R2956), .clock(clock), .in1(R2955));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3157 (.out1(R3158), .clock(clock), .in1(R3157));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3404 (.out1(R3405), .clock(clock), .in1(R3404));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3596 (.out1(R3597), .clock(clock), .in1(R3596));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3784 (.out1(R3785), .clock(clock), .in1(R3784));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4017 (.out1(R4018), .clock(clock), .in1(R4017));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4195 (.out1(R4196), .clock(clock), .in1(R4195));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4369 (.out1(R4370), .clock(clock), .in1(R4369));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4588 (.out1(R4589), .clock(clock), .in1(R4588));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4752 (.out1(R4753), .clock(clock), .in1(R4752));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4912 (.out1(R4913), .clock(clock), .in1(R4912));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5117 (.out1(R5118), .clock(clock), .in1(R5117));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5267 (.out1(R5268), .clock(clock), .in1(R5267));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5413 (.out1(R5414), .clock(clock), .in1(R5413));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5604 (.out1(R5605), .clock(clock), .in1(R5604));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5740 (.out1(R5741), .clock(clock), .in1(R5740));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5872 (.out1(R5873), .clock(clock), .in1(R5872));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6033 (.out1(R6034), .clock(clock), .in1(_455));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6034 (.out1(R6035), .clock(clock), .in1(_516));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6035 (.out1(R6036), .clock(clock), .in1(_498));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6036 (.out1(R6037), .clock(clock), .in1(_491));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6037 (.out1(R6038), .clock(clock), .in1(_480));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6038 (.out1(R6039), .clock(clock), .in1(_473));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6039 (.out1(R6040), .clock(clock), .in1(_463));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6040 (.out1(R6041), .clock(clock), .in1(_456));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op476 (.out1(_448), .in1(R5605));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op527 (.out1(_499), .in1(R6036), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op545 (.out1(_517), .in1(R6035), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op528 (.out1(_500), .in1(R6037), .in2(_499));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op509 (.out1(_481), .in1(R6038), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op492 (.out1(_464), .in1(R6040), .in2(1 'd 1));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op510 (.out1(_482), .in1(R6039), .in2(_481));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op485 (.out1(_457), .in1(R6034), .in2(R6041));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op477 (.out1(_449), .in1(_448), .in2(2 'd 2));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op546 (.out1(_518), .in1(_517), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op529 (.out1(_501), .in1(_500), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op493 (.out1(_465), .in1(_464), .in2(63 'd 6148914691236517205));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op547 (.out1(_519), .in1(_501), .in2(_518));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op511 (.out1(_483), .in1(_482), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op494 (.out1(_466), .in1(_457), .in2(_465));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2750 (.out1(R2751), .clock(clock), .in1(R2750));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2956 (.out1(R2957), .clock(clock), .in1(R2956));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3158 (.out1(R3159), .clock(clock), .in1(R3158));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3405 (.out1(R3406), .clock(clock), .in1(R3405));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3597 (.out1(R3598), .clock(clock), .in1(R3597));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3785 (.out1(R3786), .clock(clock), .in1(R3785));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4018 (.out1(R4019), .clock(clock), .in1(R4018));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4196 (.out1(R4197), .clock(clock), .in1(R4196));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4370 (.out1(R4371), .clock(clock), .in1(R4370));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4589 (.out1(R4590), .clock(clock), .in1(R4589));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4753 (.out1(R4754), .clock(clock), .in1(R4753));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4913 (.out1(R4914), .clock(clock), .in1(R4913));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5118 (.out1(R5119), .clock(clock), .in1(R5118));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5268 (.out1(R5269), .clock(clock), .in1(R5268));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5414 (.out1(R5415), .clock(clock), .in1(R5414));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5605 (.out1(R5606), .clock(clock), .in1(R5605));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5741 (.out1(R5742), .clock(clock), .in1(R5741));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5873 (.out1(R5874), .clock(clock), .in1(R5873));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6041 (.out1(R6042), .clock(clock), .in1(_449));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6042 (.out1(R6043), .clock(clock), .in1(_519));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6043 (.out1(R6044), .clock(clock), .in1(_483));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6044 (.out1(R6045), .clock(clock), .in1(_466));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op512 (.out1(_484), .in1(R6044), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op495 (.out1(_467), .in1(R6045), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op548 (.out1(_520), .in1(R6043), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op513 (.out1(_485), .in1(_467), .in2(_484));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op478 (.out1(_450), .in1(c56_popcnt_2583_D), .in2(R6042));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op549 (.out1(_521), .in1(_485), .in2(_520));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op550 (.out1(_522), .in1(_521), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2751 (.out1(R2752), .clock(clock), .in1(R2751));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2957 (.out1(R2958), .clock(clock), .in1(R2957));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3159 (.out1(R3160), .clock(clock), .in1(R3159));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3406 (.out1(R3407), .clock(clock), .in1(R3406));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3598 (.out1(R3599), .clock(clock), .in1(R3598));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3786 (.out1(R3787), .clock(clock), .in1(R3786));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4019 (.out1(R4020), .clock(clock), .in1(R4019));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4197 (.out1(R4198), .clock(clock), .in1(R4197));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4371 (.out1(R4372), .clock(clock), .in1(R4371));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4590 (.out1(R4591), .clock(clock), .in1(R4590));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4754 (.out1(R4755), .clock(clock), .in1(R4754));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4914 (.out1(R4915), .clock(clock), .in1(R4914));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5119 (.out1(R5120), .clock(clock), .in1(R5119));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5269 (.out1(R5270), .clock(clock), .in1(R5269));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5415 (.out1(R5416), .clock(clock), .in1(R5415));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5606 (.out1(R5607), .clock(clock), .in1(R5606));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5742 (.out1(R5743), .clock(clock), .in1(R5742));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5874 (.out1(R5875), .clock(clock), .in1(R5874));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6045 (.out1(R6046), .clock(clock), .in1(_450));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6046 (.out1(R6047), .clock(clock), .in1(_522));
  SRAM op479 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_451),.ADR(R6046));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op551 (.out1(_523), .in1(R6047), .in2(57 'd 72340172838076673));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2752 (.out1(R2753), .clock(clock), .in1(R2752));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2958 (.out1(R2959), .clock(clock), .in1(R2958));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3160 (.out1(R3161), .clock(clock), .in1(R3160));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3407 (.out1(R3408), .clock(clock), .in1(R3407));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3599 (.out1(R3600), .clock(clock), .in1(R3599));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3787 (.out1(R3788), .clock(clock), .in1(R3787));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4020 (.out1(R4021), .clock(clock), .in1(R4020));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4198 (.out1(R4199), .clock(clock), .in1(R4198));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4372 (.out1(R4373), .clock(clock), .in1(R4372));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4591 (.out1(R4592), .clock(clock), .in1(R4591));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4755 (.out1(R4756), .clock(clock), .in1(R4755));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4915 (.out1(R4916), .clock(clock), .in1(R4915));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5120 (.out1(R5121), .clock(clock), .in1(R5120));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5270 (.out1(R5271), .clock(clock), .in1(R5270));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5416 (.out1(R5417), .clock(clock), .in1(R5416));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5607 (.out1(R5608), .clock(clock), .in1(R5607));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5743 (.out1(R5744), .clock(clock), .in1(R5743));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5875 (.out1(R5876), .clock(clock), .in1(R5875));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6047 (.out1(R6048), .clock(clock), .in1(_451));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6048 (.out1(R6049), .clock(clock), .in1(_523));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op552 (.out1(_524), .in1(R6049), .in2(6 'd 56));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op553 (.out1(_525), .in1(_524));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op554 (.out1(ck_idx_2584), .in1(R6048), .in2(_525));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2753 (.out1(R2754), .clock(clock), .in1(R2753));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2959 (.out1(R2960), .clock(clock), .in1(R2959));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3161 (.out1(R3162), .clock(clock), .in1(R3161));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3408 (.out1(R3409), .clock(clock), .in1(R3408));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3600 (.out1(R3601), .clock(clock), .in1(R3600));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3788 (.out1(R3789), .clock(clock), .in1(R3788));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4021 (.out1(R4022), .clock(clock), .in1(R4021));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4199 (.out1(R4200), .clock(clock), .in1(R4199));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4373 (.out1(R4374), .clock(clock), .in1(R4373));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4592 (.out1(R4593), .clock(clock), .in1(R4592));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4756 (.out1(R4757), .clock(clock), .in1(R4756));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4916 (.out1(R4917), .clock(clock), .in1(R4916));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5121 (.out1(R5122), .clock(clock), .in1(R5121));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5271 (.out1(R5272), .clock(clock), .in1(R5271));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5417 (.out1(R5418), .clock(clock), .in1(R5417));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5608 (.out1(R5609), .clock(clock), .in1(R5608));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5744 (.out1(R5745), .clock(clock), .in1(R5744));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5876 (.out1(R5877), .clock(clock), .in1(R5876));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6049 (.out1(R6050), .clock(clock), .in1(ck_idx_2584));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(4), .BITSIZE_out1(32), .PRECISION(32)) op555 (.out1(_526), .in1(R6050), .in2(4 'd 8));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2754 (.out1(R2755), .clock(clock), .in1(R2754));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2960 (.out1(R2961), .clock(clock), .in1(R2960));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3162 (.out1(R3163), .clock(clock), .in1(R3162));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3409 (.out1(R3410), .clock(clock), .in1(R3409));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3601 (.out1(R3602), .clock(clock), .in1(R3601));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3789 (.out1(R3790), .clock(clock), .in1(R3789));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4022 (.out1(R4023), .clock(clock), .in1(R4022));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4200 (.out1(R4201), .clock(clock), .in1(R4200));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4374 (.out1(R4375), .clock(clock), .in1(R4374));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4593 (.out1(R4594), .clock(clock), .in1(R4593));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4757 (.out1(R4758), .clock(clock), .in1(R4757));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4917 (.out1(R4918), .clock(clock), .in1(R4917));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5122 (.out1(R5123), .clock(clock), .in1(R5122));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5272 (.out1(R5273), .clock(clock), .in1(R5272));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5418 (.out1(R5419), .clock(clock), .in1(R5418));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5609 (.out1(R5610), .clock(clock), .in1(R5609));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5745 (.out1(R5746), .clock(clock), .in1(R5745));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5877 (.out1(R5878), .clock(clock), .in1(R5877));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6050 (.out1(R6051), .clock(clock), .in1(_526));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op556 (.out1(_527), .in1(ip1_2522_D));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(8), .BITSIZE_out1(32)) op557 (.out1(_528), .in1(_527), .in2(8 'd 255));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op558 (.out1(idx_sail_2585), .in1(R6051), .in2(_528));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(3), .BITSIZE_out1(32), .PRECISION(32)) op559 (.out1(idx_2586), .in1(idx_sail_2585), .in2(3 'd 6));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2755 (.out1(R2756), .clock(clock), .in1(R2755));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2961 (.out1(R2962), .clock(clock), .in1(R2961));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3163 (.out1(R3164), .clock(clock), .in1(R3163));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3410 (.out1(R3411), .clock(clock), .in1(R3410));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3602 (.out1(R3603), .clock(clock), .in1(R3602));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3790 (.out1(R3791), .clock(clock), .in1(R3790));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4023 (.out1(R4024), .clock(clock), .in1(R4023));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4201 (.out1(R4202), .clock(clock), .in1(R4201));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4375 (.out1(R4376), .clock(clock), .in1(R4375));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4594 (.out1(R4595), .clock(clock), .in1(R4594));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4758 (.out1(R4759), .clock(clock), .in1(R4758));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4918 (.out1(R4919), .clock(clock), .in1(R4918));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5123 (.out1(R5124), .clock(clock), .in1(R5123));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5273 (.out1(R5274), .clock(clock), .in1(R5273));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5419 (.out1(R5420), .clock(clock), .in1(R5419));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5610 (.out1(R5611), .clock(clock), .in1(R5610));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5746 (.out1(R5747), .clock(clock), .in1(R5746));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5878 (.out1(R5879), .clock(clock), .in1(R5878));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6051 (.out1(R6052), .clock(clock), .in1(idx_sail_2585));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6054 (.out1(R6055), .clock(clock), .in1(idx_2586));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op561 (.out1(_529), .in1(R6055));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op562 (.out1(_530), .in1(_529), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2756 (.out1(R2757), .clock(clock), .in1(R2756));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2962 (.out1(R2963), .clock(clock), .in1(R2962));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3164 (.out1(R3165), .clock(clock), .in1(R3164));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3411 (.out1(R3412), .clock(clock), .in1(R3411));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3603 (.out1(R3604), .clock(clock), .in1(R3603));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3791 (.out1(R3792), .clock(clock), .in1(R3791));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4024 (.out1(R4025), .clock(clock), .in1(R4024));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4202 (.out1(R4203), .clock(clock), .in1(R4202));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4376 (.out1(R4377), .clock(clock), .in1(R4376));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4595 (.out1(R4596), .clock(clock), .in1(R4595));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4759 (.out1(R4760), .clock(clock), .in1(R4759));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4919 (.out1(R4920), .clock(clock), .in1(R4919));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5124 (.out1(R5125), .clock(clock), .in1(R5124));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5274 (.out1(R5275), .clock(clock), .in1(R5274));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5420 (.out1(R5421), .clock(clock), .in1(R5420));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5611 (.out1(R5612), .clock(clock), .in1(R5611));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5747 (.out1(R5748), .clock(clock), .in1(R5747));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5879 (.out1(R5880), .clock(clock), .in1(R5879));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6052 (.out1(R6053), .clock(clock), .in1(R6052));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6055 (.out1(R6056), .clock(clock), .in1(R6055));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6175 (.out1(R6176), .clock(clock), .in1(_530));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op563 (.out1(_531), .in1(c64_bitmap_2588_D), .in2(R6176));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2757 (.out1(R2758), .clock(clock), .in1(R2757));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2963 (.out1(R2964), .clock(clock), .in1(R2963));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3165 (.out1(R3166), .clock(clock), .in1(R3165));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3412 (.out1(R3413), .clock(clock), .in1(R3412));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3604 (.out1(R3605), .clock(clock), .in1(R3604));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3792 (.out1(R3793), .clock(clock), .in1(R3792));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4025 (.out1(R4026), .clock(clock), .in1(R4025));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4203 (.out1(R4204), .clock(clock), .in1(R4203));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4377 (.out1(R4378), .clock(clock), .in1(R4377));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4596 (.out1(R4597), .clock(clock), .in1(R4596));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4760 (.out1(R4761), .clock(clock), .in1(R4760));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4920 (.out1(R4921), .clock(clock), .in1(R4920));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5125 (.out1(R5126), .clock(clock), .in1(R5125));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5275 (.out1(R5276), .clock(clock), .in1(R5275));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5421 (.out1(R5422), .clock(clock), .in1(R5421));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5612 (.out1(R5613), .clock(clock), .in1(R5612));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5748 (.out1(R5749), .clock(clock), .in1(R5748));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5880 (.out1(R5881), .clock(clock), .in1(R5880));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6053 (.out1(R6054), .clock(clock), .in1(R6053));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6056 (.out1(R6057), .clock(clock), .in1(R6056));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6176 (.out1(R6177), .clock(clock), .in1(_531));
  SRAM op564 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_532),.ADR(R6177));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op560 (.out1(off_2587), .in1(R6054), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op565 (.out1(_533), .in1(64 'd 9223372036854775808), .in2(off_2587));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2758 (.out1(R2759), .clock(clock), .in1(R2758));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2964 (.out1(R2965), .clock(clock), .in1(R2964));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3166 (.out1(R3167), .clock(clock), .in1(R3166));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3413 (.out1(R3414), .clock(clock), .in1(R3413));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3605 (.out1(R3606), .clock(clock), .in1(R3605));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3793 (.out1(R3794), .clock(clock), .in1(R3793));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4026 (.out1(R4027), .clock(clock), .in1(R4026));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4204 (.out1(R4205), .clock(clock), .in1(R4204));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4378 (.out1(R4379), .clock(clock), .in1(R4378));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4597 (.out1(R4598), .clock(clock), .in1(R4597));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4761 (.out1(R4762), .clock(clock), .in1(R4761));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4921 (.out1(R4922), .clock(clock), .in1(R4921));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5126 (.out1(R5127), .clock(clock), .in1(R5126));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5276 (.out1(R5277), .clock(clock), .in1(R5276));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5422 (.out1(R5423), .clock(clock), .in1(R5422));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5613 (.out1(R5614), .clock(clock), .in1(R5613));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5749 (.out1(R5750), .clock(clock), .in1(R5749));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5881 (.out1(R5882), .clock(clock), .in1(R5881));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6057 (.out1(R6058), .clock(clock), .in1(R6057));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6177 (.out1(R6178), .clock(clock), .in1(_532));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6178 (.out1(R6179), .clock(clock), .in1(off_2587));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6295 (.out1(R6296), .clock(clock), .in1(_533));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op566 (.out1(_534), .in1(R6178), .in2(R6296));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op567 (.out1(ifout567), .in1(_534), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op628 (.out1(_595), .in1(R6058));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op629 (.out1(_596), .in1(_595), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2759 (.out1(R2760), .clock(clock), .in1(R2759));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2965 (.out1(R2966), .clock(clock), .in1(R2965));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3167 (.out1(R3168), .clock(clock), .in1(R3167));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3414 (.out1(R3415), .clock(clock), .in1(R3414));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3606 (.out1(R3607), .clock(clock), .in1(R3606));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3794 (.out1(R3795), .clock(clock), .in1(R3794));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4027 (.out1(R4028), .clock(clock), .in1(R4027));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4205 (.out1(R4206), .clock(clock), .in1(R4205));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4379 (.out1(R4380), .clock(clock), .in1(R4379));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4598 (.out1(R4599), .clock(clock), .in1(R4598));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4762 (.out1(R4763), .clock(clock), .in1(R4762));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4922 (.out1(R4923), .clock(clock), .in1(R4922));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5127 (.out1(R5128), .clock(clock), .in1(R5127));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5277 (.out1(R5278), .clock(clock), .in1(R5277));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5423 (.out1(R5424), .clock(clock), .in1(R5423));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5614 (.out1(R5615), .clock(clock), .in1(R5614));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5750 (.out1(R5751), .clock(clock), .in1(R5750));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5882 (.out1(R5883), .clock(clock), .in1(R5882));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6058 (.out1(R6059), .clock(clock), .in1(R6058));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6179 (.out1(R6180), .clock(clock), .in1(R6179));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6296 (.out1(R6297), .clock(clock), .in1(ifout567));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6420 (.out1(R6421), .clock(clock), .in1(_596));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op622 (.out1(_589), .in1(R6059));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op612 (.out1(_579), .in1(R6059));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op606 (.out1(_573), .in1(R6059));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op594 (.out1(_561), .in1(R6059));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op588 (.out1(_555), .in1(R6059));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op578 (.out1(_545), .in1(R6059));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op623 (.out1(_590), .in1(_589), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op613 (.out1(_580), .in1(_579), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op607 (.out1(_574), .in1(_573), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op595 (.out1(_562), .in1(_561), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op589 (.out1(_556), .in1(_555), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op579 (.out1(_546), .in1(_545), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op630 (.out1(_597), .in1(c64_bitmap_2588_D), .in2(R6421));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2760 (.out1(R2761), .clock(clock), .in1(R2760));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2966 (.out1(R2967), .clock(clock), .in1(R2966));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3168 (.out1(R3169), .clock(clock), .in1(R3168));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3415 (.out1(R3416), .clock(clock), .in1(R3415));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3607 (.out1(R3608), .clock(clock), .in1(R3607));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3795 (.out1(R3796), .clock(clock), .in1(R3795));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4028 (.out1(R4029), .clock(clock), .in1(R4028));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4206 (.out1(R4207), .clock(clock), .in1(R4206));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4380 (.out1(R4381), .clock(clock), .in1(R4380));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4599 (.out1(R4600), .clock(clock), .in1(R4599));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4763 (.out1(R4764), .clock(clock), .in1(R4763));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4923 (.out1(R4924), .clock(clock), .in1(R4923));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5128 (.out1(R5129), .clock(clock), .in1(R5128));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5278 (.out1(R5279), .clock(clock), .in1(R5278));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5424 (.out1(R5425), .clock(clock), .in1(R5424));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5615 (.out1(R5616), .clock(clock), .in1(R5615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5751 (.out1(R5752), .clock(clock), .in1(R5751));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5883 (.out1(R5884), .clock(clock), .in1(R5883));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6059 (.out1(R6060), .clock(clock), .in1(R6059));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6180 (.out1(R6181), .clock(clock), .in1(R6180));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6297 (.out1(R6298), .clock(clock), .in1(R6297));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6421 (.out1(R6422), .clock(clock), .in1(_590));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6422 (.out1(R6423), .clock(clock), .in1(_580));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6423 (.out1(R6424), .clock(clock), .in1(_574));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6424 (.out1(R6425), .clock(clock), .in1(_562));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6425 (.out1(R6426), .clock(clock), .in1(_556));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6426 (.out1(R6427), .clock(clock), .in1(_546));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6427 (.out1(R6428), .clock(clock), .in1(_597));
  SRAM op631 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_598),.ADR(R6428));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op572 (.out1(_539), .in1(R6060));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op573 (.out1(_540), .in1(_539), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op624 (.out1(_591), .in1(c64_bitmap_2588_D), .in2(R6422));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op614 (.out1(_581), .in1(c64_bitmap_2588_D), .in2(R6423));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op608 (.out1(_575), .in1(c64_bitmap_2588_D), .in2(R6424));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op596 (.out1(_563), .in1(c64_bitmap_2588_D), .in2(R6425));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op590 (.out1(_557), .in1(c64_bitmap_2588_D), .in2(R6426));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op580 (.out1(_547), .in1(c64_bitmap_2588_D), .in2(R6427));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2761 (.out1(R2762), .clock(clock), .in1(R2761));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2967 (.out1(R2968), .clock(clock), .in1(R2967));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3169 (.out1(R3170), .clock(clock), .in1(R3169));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3416 (.out1(R3417), .clock(clock), .in1(R3416));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3608 (.out1(R3609), .clock(clock), .in1(R3608));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3796 (.out1(R3797), .clock(clock), .in1(R3796));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4029 (.out1(R4030), .clock(clock), .in1(R4029));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4207 (.out1(R4208), .clock(clock), .in1(R4207));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4381 (.out1(R4382), .clock(clock), .in1(R4381));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4600 (.out1(R4601), .clock(clock), .in1(R4600));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4764 (.out1(R4765), .clock(clock), .in1(R4764));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4924 (.out1(R4925), .clock(clock), .in1(R4924));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5129 (.out1(R5130), .clock(clock), .in1(R5129));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5279 (.out1(R5280), .clock(clock), .in1(R5279));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5425 (.out1(R5426), .clock(clock), .in1(R5425));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5616 (.out1(R5617), .clock(clock), .in1(R5616));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5752 (.out1(R5753), .clock(clock), .in1(R5752));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5884 (.out1(R5885), .clock(clock), .in1(R5884));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6060 (.out1(R6061), .clock(clock), .in1(R6060));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6181 (.out1(R6182), .clock(clock), .in1(R6181));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6298 (.out1(R6299), .clock(clock), .in1(R6298));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6428 (.out1(R6429), .clock(clock), .in1(_598));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6429 (.out1(R6430), .clock(clock), .in1(_540));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6430 (.out1(R6431), .clock(clock), .in1(_591));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6431 (.out1(R6432), .clock(clock), .in1(_581));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6432 (.out1(R6433), .clock(clock), .in1(_575));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6433 (.out1(R6434), .clock(clock), .in1(_563));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6434 (.out1(R6435), .clock(clock), .in1(_557));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6435 (.out1(R6436), .clock(clock), .in1(_547));
  SRAM op625 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_592),.ADR(R6431));
  SRAM op615 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_582),.ADR(R6432));
  SRAM op609 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_576),.ADR(R6433));
  SRAM op597 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_564),.ADR(R6434));
  SRAM op591 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_558),.ADR(R6435));
  SRAM op581 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_548),.ADR(R6436));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op632 (.out1(_599), .in1(7 'd 64), .in2(R6182));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op574 (.out1(_541), .in1(c64_bitmap_2588_D), .in2(R6430));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op633 (.out1(_600), .in1(R6429), .in2(_599));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op626 (.out1(_593), .in1(7 'd 64), .in2(R6182));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op616 (.out1(_583), .in1(7 'd 64), .in2(R6182));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op598 (.out1(_565), .in1(7 'd 64), .in2(R6182));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2762 (.out1(R2763), .clock(clock), .in1(R2762));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2968 (.out1(R2969), .clock(clock), .in1(R2968));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3170 (.out1(R3171), .clock(clock), .in1(R3170));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3417 (.out1(R3418), .clock(clock), .in1(R3417));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3609 (.out1(R3610), .clock(clock), .in1(R3609));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3797 (.out1(R3798), .clock(clock), .in1(R3797));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4030 (.out1(R4031), .clock(clock), .in1(R4030));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4208 (.out1(R4209), .clock(clock), .in1(R4208));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4382 (.out1(R4383), .clock(clock), .in1(R4382));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4601 (.out1(R4602), .clock(clock), .in1(R4601));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4765 (.out1(R4766), .clock(clock), .in1(R4765));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4925 (.out1(R4926), .clock(clock), .in1(R4925));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5130 (.out1(R5131), .clock(clock), .in1(R5130));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5280 (.out1(R5281), .clock(clock), .in1(R5280));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5426 (.out1(R5427), .clock(clock), .in1(R5426));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5617 (.out1(R5618), .clock(clock), .in1(R5617));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5753 (.out1(R5754), .clock(clock), .in1(R5753));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5885 (.out1(R5886), .clock(clock), .in1(R5885));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6061 (.out1(R6062), .clock(clock), .in1(R6061));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6182 (.out1(R6183), .clock(clock), .in1(R6182));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6299 (.out1(R6300), .clock(clock), .in1(R6299));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6436 (.out1(R6437), .clock(clock), .in1(_592));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6437 (.out1(R6438), .clock(clock), .in1(_582));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6438 (.out1(R6439), .clock(clock), .in1(_576));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6439 (.out1(R6440), .clock(clock), .in1(_564));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6440 (.out1(R6441), .clock(clock), .in1(_558));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6441 (.out1(R6442), .clock(clock), .in1(_548));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6442 (.out1(R6443), .clock(clock), .in1(_541));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6443 (.out1(R6444), .clock(clock), .in1(_600));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6444 (.out1(R6445), .clock(clock), .in1(_593));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6445 (.out1(R6446), .clock(clock), .in1(_583));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6446 (.out1(R6447), .clock(clock), .in1(_565));
  SRAM op575 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_542),.ADR(R6443));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op634 (.out1(_601), .in1(R6444), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op627 (.out1(_594), .in1(R6437), .in2(R6445));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op617 (.out1(_584), .in1(R6438), .in2(R6446));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op610 (.out1(_577), .in1(7 'd 64), .in2(R6183));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op599 (.out1(_566), .in1(R6440), .in2(R6447));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op592 (.out1(_559), .in1(7 'd 64), .in2(R6183));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op582 (.out1(_549), .in1(7 'd 64), .in2(R6183));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op635 (.out1(_602), .in1(_601), .in2(63 'd 6148914691236517205));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op636 (.out1(_603), .in1(_594), .in2(_602));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op618 (.out1(_585), .in1(_584), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op611 (.out1(_578), .in1(R6439), .in2(_577));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op600 (.out1(_567), .in1(_566), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op593 (.out1(_560), .in1(R6441), .in2(_559));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op583 (.out1(_550), .in1(R6442), .in2(_549));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op576 (.out1(_543), .in1(7 'd 64), .in2(R6183));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2763 (.out1(R2764), .clock(clock), .in1(R2763));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2969 (.out1(R2970), .clock(clock), .in1(R2969));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3171 (.out1(R3172), .clock(clock), .in1(R3171));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3418 (.out1(R3419), .clock(clock), .in1(R3418));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3610 (.out1(R3611), .clock(clock), .in1(R3610));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3798 (.out1(R3799), .clock(clock), .in1(R3798));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4031 (.out1(R4032), .clock(clock), .in1(R4031));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4209 (.out1(R4210), .clock(clock), .in1(R4209));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4383 (.out1(R4384), .clock(clock), .in1(R4383));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4602 (.out1(R4603), .clock(clock), .in1(R4602));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4766 (.out1(R4767), .clock(clock), .in1(R4766));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4926 (.out1(R4927), .clock(clock), .in1(R4926));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5131 (.out1(R5132), .clock(clock), .in1(R5131));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5281 (.out1(R5282), .clock(clock), .in1(R5281));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5427 (.out1(R5428), .clock(clock), .in1(R5427));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5618 (.out1(R5619), .clock(clock), .in1(R5618));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5754 (.out1(R5755), .clock(clock), .in1(R5754));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5886 (.out1(R5887), .clock(clock), .in1(R5886));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6062 (.out1(R6063), .clock(clock), .in1(R6062));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6183 (.out1(R6184), .clock(clock), .in1(R6183));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6300 (.out1(R6301), .clock(clock), .in1(R6300));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6447 (.out1(R6448), .clock(clock), .in1(_542));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6448 (.out1(R6449), .clock(clock), .in1(_603));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6449 (.out1(R6450), .clock(clock), .in1(_585));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6450 (.out1(R6451), .clock(clock), .in1(_578));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6451 (.out1(R6452), .clock(clock), .in1(_567));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6452 (.out1(R6453), .clock(clock), .in1(_560));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6453 (.out1(R6454), .clock(clock), .in1(_550));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6454 (.out1(R6455), .clock(clock), .in1(_543));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op568 (.out1(_535), .in1(R6063));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op619 (.out1(_586), .in1(R6450), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op637 (.out1(_604), .in1(R6449), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op620 (.out1(_587), .in1(R6451), .in2(_586));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op601 (.out1(_568), .in1(R6452), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op584 (.out1(_551), .in1(R6454), .in2(1 'd 1));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op602 (.out1(_569), .in1(R6453), .in2(_568));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op577 (.out1(_544), .in1(R6448), .in2(R6455));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op569 (.out1(_536), .in1(_535), .in2(2 'd 2));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op638 (.out1(_605), .in1(_604), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op621 (.out1(_588), .in1(_587), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op585 (.out1(_552), .in1(_551), .in2(63 'd 6148914691236517205));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op639 (.out1(_606), .in1(_588), .in2(_605));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op603 (.out1(_570), .in1(_569), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op586 (.out1(_553), .in1(_544), .in2(_552));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2764 (.out1(R2765), .clock(clock), .in1(R2764));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2970 (.out1(R2971), .clock(clock), .in1(R2970));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3172 (.out1(R3173), .clock(clock), .in1(R3172));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3419 (.out1(R3420), .clock(clock), .in1(R3419));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3611 (.out1(R3612), .clock(clock), .in1(R3611));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3799 (.out1(R3800), .clock(clock), .in1(R3799));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4032 (.out1(R4033), .clock(clock), .in1(R4032));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4210 (.out1(R4211), .clock(clock), .in1(R4210));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4384 (.out1(R4385), .clock(clock), .in1(R4384));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4603 (.out1(R4604), .clock(clock), .in1(R4603));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4767 (.out1(R4768), .clock(clock), .in1(R4767));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4927 (.out1(R4928), .clock(clock), .in1(R4927));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5132 (.out1(R5133), .clock(clock), .in1(R5132));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5282 (.out1(R5283), .clock(clock), .in1(R5282));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5428 (.out1(R5429), .clock(clock), .in1(R5428));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5619 (.out1(R5620), .clock(clock), .in1(R5619));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5755 (.out1(R5756), .clock(clock), .in1(R5755));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5887 (.out1(R5888), .clock(clock), .in1(R5887));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6063 (.out1(R6064), .clock(clock), .in1(R6063));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6184 (.out1(R6185), .clock(clock), .in1(R6184));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6301 (.out1(R6302), .clock(clock), .in1(R6301));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6455 (.out1(R6456), .clock(clock), .in1(_536));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6456 (.out1(R6457), .clock(clock), .in1(_606));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6457 (.out1(R6458), .clock(clock), .in1(_570));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6458 (.out1(R6459), .clock(clock), .in1(_553));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op604 (.out1(_571), .in1(R6458), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op587 (.out1(_554), .in1(R6459), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op640 (.out1(_607), .in1(R6457), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op605 (.out1(_572), .in1(_554), .in2(_571));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op570 (.out1(_537), .in1(c64_popcnt_2593_D), .in2(R6456));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op641 (.out1(_608), .in1(_572), .in2(_607));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op642 (.out1(_609), .in1(_608), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2765 (.out1(R2766), .clock(clock), .in1(R2765));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2971 (.out1(R2972), .clock(clock), .in1(R2971));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3173 (.out1(R3174), .clock(clock), .in1(R3173));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3420 (.out1(R3421), .clock(clock), .in1(R3420));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3612 (.out1(R3613), .clock(clock), .in1(R3612));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3800 (.out1(R3801), .clock(clock), .in1(R3800));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4033 (.out1(R4034), .clock(clock), .in1(R4033));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4211 (.out1(R4212), .clock(clock), .in1(R4211));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4385 (.out1(R4386), .clock(clock), .in1(R4385));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4604 (.out1(R4605), .clock(clock), .in1(R4604));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4768 (.out1(R4769), .clock(clock), .in1(R4768));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4928 (.out1(R4929), .clock(clock), .in1(R4928));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5133 (.out1(R5134), .clock(clock), .in1(R5133));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5283 (.out1(R5284), .clock(clock), .in1(R5283));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5429 (.out1(R5430), .clock(clock), .in1(R5429));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5620 (.out1(R5621), .clock(clock), .in1(R5620));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5756 (.out1(R5757), .clock(clock), .in1(R5756));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5888 (.out1(R5889), .clock(clock), .in1(R5888));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6064 (.out1(R6065), .clock(clock), .in1(R6064));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6185 (.out1(R6186), .clock(clock), .in1(R6185));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6302 (.out1(R6303), .clock(clock), .in1(R6302));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6459 (.out1(R6460), .clock(clock), .in1(_537));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6460 (.out1(R6461), .clock(clock), .in1(_609));
  SRAM op571 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_538),.ADR(R6460));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op643 (.out1(_610), .in1(R6461), .in2(57 'd 72340172838076673));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2766 (.out1(R2767), .clock(clock), .in1(R2766));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2972 (.out1(R2973), .clock(clock), .in1(R2972));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3174 (.out1(R3175), .clock(clock), .in1(R3174));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3421 (.out1(R3422), .clock(clock), .in1(R3421));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3613 (.out1(R3614), .clock(clock), .in1(R3613));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3801 (.out1(R3802), .clock(clock), .in1(R3801));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4034 (.out1(R4035), .clock(clock), .in1(R4034));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4212 (.out1(R4213), .clock(clock), .in1(R4212));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4386 (.out1(R4387), .clock(clock), .in1(R4386));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4605 (.out1(R4606), .clock(clock), .in1(R4605));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4769 (.out1(R4770), .clock(clock), .in1(R4769));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4929 (.out1(R4930), .clock(clock), .in1(R4929));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5134 (.out1(R5135), .clock(clock), .in1(R5134));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5284 (.out1(R5285), .clock(clock), .in1(R5284));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5430 (.out1(R5431), .clock(clock), .in1(R5430));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5621 (.out1(R5622), .clock(clock), .in1(R5621));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5757 (.out1(R5758), .clock(clock), .in1(R5757));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5889 (.out1(R5890), .clock(clock), .in1(R5889));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6065 (.out1(R6066), .clock(clock), .in1(R6065));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6186 (.out1(R6187), .clock(clock), .in1(R6186));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6303 (.out1(R6304), .clock(clock), .in1(R6303));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6461 (.out1(R6462), .clock(clock), .in1(_538));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6462 (.out1(R6463), .clock(clock), .in1(_610));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op644 (.out1(_611), .in1(R6463), .in2(6 'd 56));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op645 (.out1(_612), .in1(_611));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op646 (.out1(ck_idx_2594), .in1(R6462), .in2(_612));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2767 (.out1(R2768), .clock(clock), .in1(R2767));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2973 (.out1(R2974), .clock(clock), .in1(R2973));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3175 (.out1(R3176), .clock(clock), .in1(R3175));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3422 (.out1(R3423), .clock(clock), .in1(R3422));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3614 (.out1(R3615), .clock(clock), .in1(R3614));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3802 (.out1(R3803), .clock(clock), .in1(R3802));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4035 (.out1(R4036), .clock(clock), .in1(R4035));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4213 (.out1(R4214), .clock(clock), .in1(R4213));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4387 (.out1(R4388), .clock(clock), .in1(R4387));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4606 (.out1(R4607), .clock(clock), .in1(R4606));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4770 (.out1(R4771), .clock(clock), .in1(R4770));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4930 (.out1(R4931), .clock(clock), .in1(R4930));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5135 (.out1(R5136), .clock(clock), .in1(R5135));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5285 (.out1(R5286), .clock(clock), .in1(R5285));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5431 (.out1(R5432), .clock(clock), .in1(R5431));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5622 (.out1(R5623), .clock(clock), .in1(R5622));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5758 (.out1(R5759), .clock(clock), .in1(R5758));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5890 (.out1(R5891), .clock(clock), .in1(R5890));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6066 (.out1(R6067), .clock(clock), .in1(R6066));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6187 (.out1(R6188), .clock(clock), .in1(R6187));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6304 (.out1(R6305), .clock(clock), .in1(R6304));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6463 (.out1(R6464), .clock(clock), .in1(ck_idx_2594));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(4), .BITSIZE_out1(32), .PRECISION(32)) op647 (.out1(_613), .in1(R6464), .in2(4 'd 8));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op648 (.out1(_614), .in1(ip2_2595_D), .in2(6 'd 56));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2768 (.out1(R2769), .clock(clock), .in1(R2768));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2974 (.out1(R2975), .clock(clock), .in1(R2974));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3176 (.out1(R3177), .clock(clock), .in1(R3176));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3423 (.out1(R3424), .clock(clock), .in1(R3423));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3615 (.out1(R3616), .clock(clock), .in1(R3615));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3803 (.out1(R3804), .clock(clock), .in1(R3803));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4036 (.out1(R4037), .clock(clock), .in1(R4036));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4214 (.out1(R4215), .clock(clock), .in1(R4214));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4388 (.out1(R4389), .clock(clock), .in1(R4388));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4607 (.out1(R4608), .clock(clock), .in1(R4607));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4771 (.out1(R4772), .clock(clock), .in1(R4771));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4931 (.out1(R4932), .clock(clock), .in1(R4931));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5136 (.out1(R5137), .clock(clock), .in1(R5136));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5286 (.out1(R5287), .clock(clock), .in1(R5286));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5432 (.out1(R5433), .clock(clock), .in1(R5432));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5623 (.out1(R5624), .clock(clock), .in1(R5623));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5759 (.out1(R5760), .clock(clock), .in1(R5759));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5891 (.out1(R5892), .clock(clock), .in1(R5891));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6067 (.out1(R6068), .clock(clock), .in1(R6067));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6188 (.out1(R6189), .clock(clock), .in1(R6188));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6305 (.out1(R6306), .clock(clock), .in1(R6305));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6464 (.out1(R6465), .clock(clock), .in1(_613));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6465 (.out1(R6466), .clock(clock), .in1(_614));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op649 (.out1(_615), .in1(R6466));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op650 (.out1(idx_sail_2596), .in1(R6465), .in2(_615));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(3), .BITSIZE_out1(32), .PRECISION(32)) op651 (.out1(idx_2597), .in1(idx_sail_2596), .in2(3 'd 6));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2769 (.out1(R2770), .clock(clock), .in1(R2769));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2975 (.out1(R2976), .clock(clock), .in1(R2975));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3177 (.out1(R3178), .clock(clock), .in1(R3177));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3424 (.out1(R3425), .clock(clock), .in1(R3424));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3616 (.out1(R3617), .clock(clock), .in1(R3616));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3804 (.out1(R3805), .clock(clock), .in1(R3804));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4037 (.out1(R4038), .clock(clock), .in1(R4037));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4215 (.out1(R4216), .clock(clock), .in1(R4215));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4389 (.out1(R4390), .clock(clock), .in1(R4389));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4608 (.out1(R4609), .clock(clock), .in1(R4608));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4772 (.out1(R4773), .clock(clock), .in1(R4772));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4932 (.out1(R4933), .clock(clock), .in1(R4932));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5137 (.out1(R5138), .clock(clock), .in1(R5137));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5287 (.out1(R5288), .clock(clock), .in1(R5287));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5433 (.out1(R5434), .clock(clock), .in1(R5433));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5624 (.out1(R5625), .clock(clock), .in1(R5624));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5760 (.out1(R5761), .clock(clock), .in1(R5760));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5892 (.out1(R5893), .clock(clock), .in1(R5892));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6068 (.out1(R6069), .clock(clock), .in1(R6068));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6189 (.out1(R6190), .clock(clock), .in1(R6189));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6306 (.out1(R6307), .clock(clock), .in1(R6306));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6466 (.out1(R6467), .clock(clock), .in1(idx_sail_2596));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6469 (.out1(R6470), .clock(clock), .in1(idx_2597));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op653 (.out1(_616), .in1(R6470));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op654 (.out1(_617), .in1(_616), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2770 (.out1(R2771), .clock(clock), .in1(R2770));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2976 (.out1(R2977), .clock(clock), .in1(R2976));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3178 (.out1(R3179), .clock(clock), .in1(R3178));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3425 (.out1(R3426), .clock(clock), .in1(R3425));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3617 (.out1(R3618), .clock(clock), .in1(R3617));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3805 (.out1(R3806), .clock(clock), .in1(R3805));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4038 (.out1(R4039), .clock(clock), .in1(R4038));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4216 (.out1(R4217), .clock(clock), .in1(R4216));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4390 (.out1(R4391), .clock(clock), .in1(R4390));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4609 (.out1(R4610), .clock(clock), .in1(R4609));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4773 (.out1(R4774), .clock(clock), .in1(R4773));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4933 (.out1(R4934), .clock(clock), .in1(R4933));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5138 (.out1(R5139), .clock(clock), .in1(R5138));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5288 (.out1(R5289), .clock(clock), .in1(R5288));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5434 (.out1(R5435), .clock(clock), .in1(R5434));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5625 (.out1(R5626), .clock(clock), .in1(R5625));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5761 (.out1(R5762), .clock(clock), .in1(R5761));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5893 (.out1(R5894), .clock(clock), .in1(R5893));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6069 (.out1(R6070), .clock(clock), .in1(R6069));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6190 (.out1(R6191), .clock(clock), .in1(R6190));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6307 (.out1(R6308), .clock(clock), .in1(R6307));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6467 (.out1(R6468), .clock(clock), .in1(R6467));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6470 (.out1(R6471), .clock(clock), .in1(R6470));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6576 (.out1(R6577), .clock(clock), .in1(_617));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op655 (.out1(_618), .in1(c72_bitmap_2599_D), .in2(R6577));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2771 (.out1(R2772), .clock(clock), .in1(R2771));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2977 (.out1(R2978), .clock(clock), .in1(R2977));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3179 (.out1(R3180), .clock(clock), .in1(R3179));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3426 (.out1(R3427), .clock(clock), .in1(R3426));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3618 (.out1(R3619), .clock(clock), .in1(R3618));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3806 (.out1(R3807), .clock(clock), .in1(R3806));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4039 (.out1(R4040), .clock(clock), .in1(R4039));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4217 (.out1(R4218), .clock(clock), .in1(R4217));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4391 (.out1(R4392), .clock(clock), .in1(R4391));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4610 (.out1(R4611), .clock(clock), .in1(R4610));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4774 (.out1(R4775), .clock(clock), .in1(R4774));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4934 (.out1(R4935), .clock(clock), .in1(R4934));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5139 (.out1(R5140), .clock(clock), .in1(R5139));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5289 (.out1(R5290), .clock(clock), .in1(R5289));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5435 (.out1(R5436), .clock(clock), .in1(R5435));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5626 (.out1(R5627), .clock(clock), .in1(R5626));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5762 (.out1(R5763), .clock(clock), .in1(R5762));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5894 (.out1(R5895), .clock(clock), .in1(R5894));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6070 (.out1(R6071), .clock(clock), .in1(R6070));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6191 (.out1(R6192), .clock(clock), .in1(R6191));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6308 (.out1(R6309), .clock(clock), .in1(R6308));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6468 (.out1(R6469), .clock(clock), .in1(R6468));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6471 (.out1(R6472), .clock(clock), .in1(R6471));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6577 (.out1(R6578), .clock(clock), .in1(_618));
  SRAM op656 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_619),.ADR(R6578));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op652 (.out1(off_2598), .in1(R6469), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op657 (.out1(_620), .in1(64 'd 9223372036854775808), .in2(off_2598));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2772 (.out1(R2773), .clock(clock), .in1(R2772));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2978 (.out1(R2979), .clock(clock), .in1(R2978));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3180 (.out1(R3181), .clock(clock), .in1(R3180));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3427 (.out1(R3428), .clock(clock), .in1(R3427));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3619 (.out1(R3620), .clock(clock), .in1(R3619));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3807 (.out1(R3808), .clock(clock), .in1(R3807));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4040 (.out1(R4041), .clock(clock), .in1(R4040));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4218 (.out1(R4219), .clock(clock), .in1(R4218));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4392 (.out1(R4393), .clock(clock), .in1(R4392));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4611 (.out1(R4612), .clock(clock), .in1(R4611));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4775 (.out1(R4776), .clock(clock), .in1(R4775));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4935 (.out1(R4936), .clock(clock), .in1(R4935));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5140 (.out1(R5141), .clock(clock), .in1(R5140));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5290 (.out1(R5291), .clock(clock), .in1(R5290));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5436 (.out1(R5437), .clock(clock), .in1(R5436));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5627 (.out1(R5628), .clock(clock), .in1(R5627));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5763 (.out1(R5764), .clock(clock), .in1(R5763));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5895 (.out1(R5896), .clock(clock), .in1(R5895));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6071 (.out1(R6072), .clock(clock), .in1(R6071));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6192 (.out1(R6193), .clock(clock), .in1(R6192));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6309 (.out1(R6310), .clock(clock), .in1(R6309));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6472 (.out1(R6473), .clock(clock), .in1(R6472));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6578 (.out1(R6579), .clock(clock), .in1(_619));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6579 (.out1(R6580), .clock(clock), .in1(off_2598));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6682 (.out1(R6683), .clock(clock), .in1(_620));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op658 (.out1(_621), .in1(R6579), .in2(R6683));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op659 (.out1(ifout659), .in1(_621), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op720 (.out1(_682), .in1(R6473));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op721 (.out1(_683), .in1(_682), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2773 (.out1(R2774), .clock(clock), .in1(R2773));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2979 (.out1(R2980), .clock(clock), .in1(R2979));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3181 (.out1(R3182), .clock(clock), .in1(R3181));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3428 (.out1(R3429), .clock(clock), .in1(R3428));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3620 (.out1(R3621), .clock(clock), .in1(R3620));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3808 (.out1(R3809), .clock(clock), .in1(R3808));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4041 (.out1(R4042), .clock(clock), .in1(R4041));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4219 (.out1(R4220), .clock(clock), .in1(R4219));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4393 (.out1(R4394), .clock(clock), .in1(R4393));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4612 (.out1(R4613), .clock(clock), .in1(R4612));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4776 (.out1(R4777), .clock(clock), .in1(R4776));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4936 (.out1(R4937), .clock(clock), .in1(R4936));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5141 (.out1(R5142), .clock(clock), .in1(R5141));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5291 (.out1(R5292), .clock(clock), .in1(R5291));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5437 (.out1(R5438), .clock(clock), .in1(R5437));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5628 (.out1(R5629), .clock(clock), .in1(R5628));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5764 (.out1(R5765), .clock(clock), .in1(R5764));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5896 (.out1(R5897), .clock(clock), .in1(R5896));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6072 (.out1(R6073), .clock(clock), .in1(R6072));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6193 (.out1(R6194), .clock(clock), .in1(R6193));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6310 (.out1(R6311), .clock(clock), .in1(R6310));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6473 (.out1(R6474), .clock(clock), .in1(R6473));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6580 (.out1(R6581), .clock(clock), .in1(R6580));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6683 (.out1(R6684), .clock(clock), .in1(ifout659));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6792 (.out1(R6793), .clock(clock), .in1(_683));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op714 (.out1(_676), .in1(R6474));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op704 (.out1(_666), .in1(R6474));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op698 (.out1(_660), .in1(R6474));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op686 (.out1(_648), .in1(R6474));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op680 (.out1(_642), .in1(R6474));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op670 (.out1(_632), .in1(R6474));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op715 (.out1(_677), .in1(_676), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op705 (.out1(_667), .in1(_666), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op699 (.out1(_661), .in1(_660), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op687 (.out1(_649), .in1(_648), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op681 (.out1(_643), .in1(_642), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op671 (.out1(_633), .in1(_632), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op722 (.out1(_684), .in1(c72_bitmap_2599_D), .in2(R6793));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2774 (.out1(R2775), .clock(clock), .in1(R2774));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2980 (.out1(R2981), .clock(clock), .in1(R2980));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3182 (.out1(R3183), .clock(clock), .in1(R3182));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3429 (.out1(R3430), .clock(clock), .in1(R3429));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3621 (.out1(R3622), .clock(clock), .in1(R3621));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3809 (.out1(R3810), .clock(clock), .in1(R3809));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4042 (.out1(R4043), .clock(clock), .in1(R4042));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4220 (.out1(R4221), .clock(clock), .in1(R4220));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4394 (.out1(R4395), .clock(clock), .in1(R4394));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4613 (.out1(R4614), .clock(clock), .in1(R4613));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4777 (.out1(R4778), .clock(clock), .in1(R4777));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4937 (.out1(R4938), .clock(clock), .in1(R4937));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5142 (.out1(R5143), .clock(clock), .in1(R5142));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5292 (.out1(R5293), .clock(clock), .in1(R5292));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5438 (.out1(R5439), .clock(clock), .in1(R5438));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5629 (.out1(R5630), .clock(clock), .in1(R5629));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5765 (.out1(R5766), .clock(clock), .in1(R5765));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5897 (.out1(R5898), .clock(clock), .in1(R5897));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6073 (.out1(R6074), .clock(clock), .in1(R6073));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6194 (.out1(R6195), .clock(clock), .in1(R6194));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6311 (.out1(R6312), .clock(clock), .in1(R6311));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6474 (.out1(R6475), .clock(clock), .in1(R6474));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6581 (.out1(R6582), .clock(clock), .in1(R6581));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6684 (.out1(R6685), .clock(clock), .in1(R6684));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6793 (.out1(R6794), .clock(clock), .in1(_677));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6794 (.out1(R6795), .clock(clock), .in1(_667));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6795 (.out1(R6796), .clock(clock), .in1(_661));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6796 (.out1(R6797), .clock(clock), .in1(_649));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6797 (.out1(R6798), .clock(clock), .in1(_643));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6798 (.out1(R6799), .clock(clock), .in1(_633));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6799 (.out1(R6800), .clock(clock), .in1(_684));
  SRAM op723 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_685),.ADR(R6800));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op664 (.out1(_626), .in1(R6475));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op665 (.out1(_627), .in1(_626), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op716 (.out1(_678), .in1(c72_bitmap_2599_D), .in2(R6794));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op706 (.out1(_668), .in1(c72_bitmap_2599_D), .in2(R6795));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op700 (.out1(_662), .in1(c72_bitmap_2599_D), .in2(R6796));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op688 (.out1(_650), .in1(c72_bitmap_2599_D), .in2(R6797));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op682 (.out1(_644), .in1(c72_bitmap_2599_D), .in2(R6798));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op672 (.out1(_634), .in1(c72_bitmap_2599_D), .in2(R6799));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2775 (.out1(R2776), .clock(clock), .in1(R2775));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2981 (.out1(R2982), .clock(clock), .in1(R2981));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3183 (.out1(R3184), .clock(clock), .in1(R3183));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3430 (.out1(R3431), .clock(clock), .in1(R3430));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3622 (.out1(R3623), .clock(clock), .in1(R3622));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3810 (.out1(R3811), .clock(clock), .in1(R3810));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4043 (.out1(R4044), .clock(clock), .in1(R4043));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4221 (.out1(R4222), .clock(clock), .in1(R4221));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4395 (.out1(R4396), .clock(clock), .in1(R4395));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4614 (.out1(R4615), .clock(clock), .in1(R4614));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4778 (.out1(R4779), .clock(clock), .in1(R4778));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4938 (.out1(R4939), .clock(clock), .in1(R4938));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5143 (.out1(R5144), .clock(clock), .in1(R5143));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5293 (.out1(R5294), .clock(clock), .in1(R5293));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5439 (.out1(R5440), .clock(clock), .in1(R5439));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5630 (.out1(R5631), .clock(clock), .in1(R5630));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5766 (.out1(R5767), .clock(clock), .in1(R5766));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5898 (.out1(R5899), .clock(clock), .in1(R5898));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6074 (.out1(R6075), .clock(clock), .in1(R6074));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6195 (.out1(R6196), .clock(clock), .in1(R6195));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6312 (.out1(R6313), .clock(clock), .in1(R6312));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6475 (.out1(R6476), .clock(clock), .in1(R6475));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6582 (.out1(R6583), .clock(clock), .in1(R6582));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6685 (.out1(R6686), .clock(clock), .in1(R6685));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6800 (.out1(R6801), .clock(clock), .in1(_685));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6801 (.out1(R6802), .clock(clock), .in1(_627));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6802 (.out1(R6803), .clock(clock), .in1(_678));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6803 (.out1(R6804), .clock(clock), .in1(_668));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6804 (.out1(R6805), .clock(clock), .in1(_662));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6805 (.out1(R6806), .clock(clock), .in1(_650));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6806 (.out1(R6807), .clock(clock), .in1(_644));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6807 (.out1(R6808), .clock(clock), .in1(_634));
  SRAM op717 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_679),.ADR(R6803));
  SRAM op707 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_669),.ADR(R6804));
  SRAM op701 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_663),.ADR(R6805));
  SRAM op689 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_651),.ADR(R6806));
  SRAM op683 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_645),.ADR(R6807));
  SRAM op673 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_635),.ADR(R6808));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op724 (.out1(_686), .in1(7 'd 64), .in2(R6583));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op666 (.out1(_628), .in1(c72_bitmap_2599_D), .in2(R6802));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op725 (.out1(_687), .in1(R6801), .in2(_686));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op718 (.out1(_680), .in1(7 'd 64), .in2(R6583));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op708 (.out1(_670), .in1(7 'd 64), .in2(R6583));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op690 (.out1(_652), .in1(7 'd 64), .in2(R6583));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2776 (.out1(R2777), .clock(clock), .in1(R2776));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2982 (.out1(R2983), .clock(clock), .in1(R2982));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3184 (.out1(R3185), .clock(clock), .in1(R3184));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3431 (.out1(R3432), .clock(clock), .in1(R3431));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3623 (.out1(R3624), .clock(clock), .in1(R3623));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3811 (.out1(R3812), .clock(clock), .in1(R3811));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4044 (.out1(R4045), .clock(clock), .in1(R4044));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4222 (.out1(R4223), .clock(clock), .in1(R4222));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4396 (.out1(R4397), .clock(clock), .in1(R4396));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4615 (.out1(R4616), .clock(clock), .in1(R4615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4779 (.out1(R4780), .clock(clock), .in1(R4779));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4939 (.out1(R4940), .clock(clock), .in1(R4939));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5144 (.out1(R5145), .clock(clock), .in1(R5144));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5294 (.out1(R5295), .clock(clock), .in1(R5294));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5440 (.out1(R5441), .clock(clock), .in1(R5440));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5631 (.out1(R5632), .clock(clock), .in1(R5631));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5767 (.out1(R5768), .clock(clock), .in1(R5767));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5899 (.out1(R5900), .clock(clock), .in1(R5899));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6075 (.out1(R6076), .clock(clock), .in1(R6075));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6196 (.out1(R6197), .clock(clock), .in1(R6196));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6313 (.out1(R6314), .clock(clock), .in1(R6313));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6476 (.out1(R6477), .clock(clock), .in1(R6476));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6583 (.out1(R6584), .clock(clock), .in1(R6583));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6686 (.out1(R6687), .clock(clock), .in1(R6686));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6808 (.out1(R6809), .clock(clock), .in1(_679));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6809 (.out1(R6810), .clock(clock), .in1(_669));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6810 (.out1(R6811), .clock(clock), .in1(_663));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6811 (.out1(R6812), .clock(clock), .in1(_651));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6812 (.out1(R6813), .clock(clock), .in1(_645));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6813 (.out1(R6814), .clock(clock), .in1(_635));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6814 (.out1(R6815), .clock(clock), .in1(_628));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6815 (.out1(R6816), .clock(clock), .in1(_687));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6816 (.out1(R6817), .clock(clock), .in1(_680));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6817 (.out1(R6818), .clock(clock), .in1(_670));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6818 (.out1(R6819), .clock(clock), .in1(_652));
  SRAM op667 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_629),.ADR(R6815));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op726 (.out1(_688), .in1(R6816), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op719 (.out1(_681), .in1(R6809), .in2(R6817));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op709 (.out1(_671), .in1(R6810), .in2(R6818));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op702 (.out1(_664), .in1(7 'd 64), .in2(R6584));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op691 (.out1(_653), .in1(R6812), .in2(R6819));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op684 (.out1(_646), .in1(7 'd 64), .in2(R6584));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op674 (.out1(_636), .in1(7 'd 64), .in2(R6584));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op727 (.out1(_689), .in1(_688), .in2(63 'd 6148914691236517205));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op728 (.out1(_690), .in1(_681), .in2(_689));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op710 (.out1(_672), .in1(_671), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op703 (.out1(_665), .in1(R6811), .in2(_664));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op692 (.out1(_654), .in1(_653), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op685 (.out1(_647), .in1(R6813), .in2(_646));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op675 (.out1(_637), .in1(R6814), .in2(_636));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op668 (.out1(_630), .in1(7 'd 64), .in2(R6584));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2777 (.out1(R2778), .clock(clock), .in1(R2777));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2983 (.out1(R2984), .clock(clock), .in1(R2983));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3185 (.out1(R3186), .clock(clock), .in1(R3185));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3432 (.out1(R3433), .clock(clock), .in1(R3432));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3624 (.out1(R3625), .clock(clock), .in1(R3624));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3812 (.out1(R3813), .clock(clock), .in1(R3812));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4045 (.out1(R4046), .clock(clock), .in1(R4045));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4223 (.out1(R4224), .clock(clock), .in1(R4223));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4397 (.out1(R4398), .clock(clock), .in1(R4397));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4616 (.out1(R4617), .clock(clock), .in1(R4616));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4780 (.out1(R4781), .clock(clock), .in1(R4780));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4940 (.out1(R4941), .clock(clock), .in1(R4940));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5145 (.out1(R5146), .clock(clock), .in1(R5145));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5295 (.out1(R5296), .clock(clock), .in1(R5295));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5441 (.out1(R5442), .clock(clock), .in1(R5441));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5632 (.out1(R5633), .clock(clock), .in1(R5632));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5768 (.out1(R5769), .clock(clock), .in1(R5768));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5900 (.out1(R5901), .clock(clock), .in1(R5900));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6076 (.out1(R6077), .clock(clock), .in1(R6076));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6197 (.out1(R6198), .clock(clock), .in1(R6197));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6314 (.out1(R6315), .clock(clock), .in1(R6314));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6477 (.out1(R6478), .clock(clock), .in1(R6477));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6584 (.out1(R6585), .clock(clock), .in1(R6584));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6687 (.out1(R6688), .clock(clock), .in1(R6687));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6819 (.out1(R6820), .clock(clock), .in1(_629));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6820 (.out1(R6821), .clock(clock), .in1(_690));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6821 (.out1(R6822), .clock(clock), .in1(_672));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6822 (.out1(R6823), .clock(clock), .in1(_665));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6823 (.out1(R6824), .clock(clock), .in1(_654));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6824 (.out1(R6825), .clock(clock), .in1(_647));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6825 (.out1(R6826), .clock(clock), .in1(_637));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6826 (.out1(R6827), .clock(clock), .in1(_630));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op660 (.out1(_622), .in1(R6478));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op711 (.out1(_673), .in1(R6822), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op729 (.out1(_691), .in1(R6821), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op712 (.out1(_674), .in1(R6823), .in2(_673));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op693 (.out1(_655), .in1(R6824), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op676 (.out1(_638), .in1(R6826), .in2(1 'd 1));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op694 (.out1(_656), .in1(R6825), .in2(_655));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op669 (.out1(_631), .in1(R6820), .in2(R6827));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op661 (.out1(_623), .in1(_622), .in2(2 'd 2));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op730 (.out1(_692), .in1(_691), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op713 (.out1(_675), .in1(_674), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op677 (.out1(_639), .in1(_638), .in2(63 'd 6148914691236517205));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op731 (.out1(_693), .in1(_675), .in2(_692));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op695 (.out1(_657), .in1(_656), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op678 (.out1(_640), .in1(_631), .in2(_639));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2778 (.out1(R2779), .clock(clock), .in1(R2778));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2984 (.out1(R2985), .clock(clock), .in1(R2984));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3186 (.out1(R3187), .clock(clock), .in1(R3186));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3433 (.out1(R3434), .clock(clock), .in1(R3433));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3625 (.out1(R3626), .clock(clock), .in1(R3625));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3813 (.out1(R3814), .clock(clock), .in1(R3813));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4046 (.out1(R4047), .clock(clock), .in1(R4046));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4224 (.out1(R4225), .clock(clock), .in1(R4224));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4398 (.out1(R4399), .clock(clock), .in1(R4398));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4617 (.out1(R4618), .clock(clock), .in1(R4617));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4781 (.out1(R4782), .clock(clock), .in1(R4781));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4941 (.out1(R4942), .clock(clock), .in1(R4941));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5146 (.out1(R5147), .clock(clock), .in1(R5146));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5296 (.out1(R5297), .clock(clock), .in1(R5296));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5442 (.out1(R5443), .clock(clock), .in1(R5442));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5633 (.out1(R5634), .clock(clock), .in1(R5633));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5769 (.out1(R5770), .clock(clock), .in1(R5769));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5901 (.out1(R5902), .clock(clock), .in1(R5901));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6077 (.out1(R6078), .clock(clock), .in1(R6077));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6198 (.out1(R6199), .clock(clock), .in1(R6198));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6315 (.out1(R6316), .clock(clock), .in1(R6315));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6478 (.out1(R6479), .clock(clock), .in1(R6478));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6585 (.out1(R6586), .clock(clock), .in1(R6585));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6688 (.out1(R6689), .clock(clock), .in1(R6688));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6827 (.out1(R6828), .clock(clock), .in1(_623));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6828 (.out1(R6829), .clock(clock), .in1(_693));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6829 (.out1(R6830), .clock(clock), .in1(_657));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6830 (.out1(R6831), .clock(clock), .in1(_640));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op696 (.out1(_658), .in1(R6830), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op679 (.out1(_641), .in1(R6831), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op732 (.out1(_694), .in1(R6829), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op697 (.out1(_659), .in1(_641), .in2(_658));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op662 (.out1(_624), .in1(c72_popcnt_2604_D), .in2(R6828));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op733 (.out1(_695), .in1(_659), .in2(_694));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op734 (.out1(_696), .in1(_695), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2779 (.out1(R2780), .clock(clock), .in1(R2779));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2985 (.out1(R2986), .clock(clock), .in1(R2985));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3187 (.out1(R3188), .clock(clock), .in1(R3187));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3434 (.out1(R3435), .clock(clock), .in1(R3434));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3626 (.out1(R3627), .clock(clock), .in1(R3626));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3814 (.out1(R3815), .clock(clock), .in1(R3814));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4047 (.out1(R4048), .clock(clock), .in1(R4047));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4225 (.out1(R4226), .clock(clock), .in1(R4225));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4399 (.out1(R4400), .clock(clock), .in1(R4399));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4618 (.out1(R4619), .clock(clock), .in1(R4618));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4782 (.out1(R4783), .clock(clock), .in1(R4782));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4942 (.out1(R4943), .clock(clock), .in1(R4942));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5147 (.out1(R5148), .clock(clock), .in1(R5147));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5297 (.out1(R5298), .clock(clock), .in1(R5297));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5443 (.out1(R5444), .clock(clock), .in1(R5443));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5634 (.out1(R5635), .clock(clock), .in1(R5634));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5770 (.out1(R5771), .clock(clock), .in1(R5770));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5902 (.out1(R5903), .clock(clock), .in1(R5902));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6078 (.out1(R6079), .clock(clock), .in1(R6078));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6199 (.out1(R6200), .clock(clock), .in1(R6199));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6316 (.out1(R6317), .clock(clock), .in1(R6316));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6479 (.out1(R6480), .clock(clock), .in1(R6479));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6586 (.out1(R6587), .clock(clock), .in1(R6586));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6689 (.out1(R6690), .clock(clock), .in1(R6689));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6831 (.out1(R6832), .clock(clock), .in1(_624));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6832 (.out1(R6833), .clock(clock), .in1(_696));
  SRAM op663 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_625),.ADR(R6832));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op735 (.out1(_697), .in1(R6833), .in2(57 'd 72340172838076673));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2780 (.out1(R2781), .clock(clock), .in1(R2780));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2986 (.out1(R2987), .clock(clock), .in1(R2986));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3188 (.out1(R3189), .clock(clock), .in1(R3188));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3435 (.out1(R3436), .clock(clock), .in1(R3435));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3627 (.out1(R3628), .clock(clock), .in1(R3627));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3815 (.out1(R3816), .clock(clock), .in1(R3815));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4048 (.out1(R4049), .clock(clock), .in1(R4048));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4226 (.out1(R4227), .clock(clock), .in1(R4226));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4400 (.out1(R4401), .clock(clock), .in1(R4400));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4619 (.out1(R4620), .clock(clock), .in1(R4619));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4783 (.out1(R4784), .clock(clock), .in1(R4783));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4943 (.out1(R4944), .clock(clock), .in1(R4943));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5148 (.out1(R5149), .clock(clock), .in1(R5148));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5298 (.out1(R5299), .clock(clock), .in1(R5298));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5444 (.out1(R5445), .clock(clock), .in1(R5444));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5635 (.out1(R5636), .clock(clock), .in1(R5635));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5771 (.out1(R5772), .clock(clock), .in1(R5771));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5903 (.out1(R5904), .clock(clock), .in1(R5903));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6079 (.out1(R6080), .clock(clock), .in1(R6079));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6200 (.out1(R6201), .clock(clock), .in1(R6200));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6317 (.out1(R6318), .clock(clock), .in1(R6317));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6480 (.out1(R6481), .clock(clock), .in1(R6480));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6587 (.out1(R6588), .clock(clock), .in1(R6587));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6690 (.out1(R6691), .clock(clock), .in1(R6690));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6833 (.out1(R6834), .clock(clock), .in1(_625));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6834 (.out1(R6835), .clock(clock), .in1(_697));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op736 (.out1(_698), .in1(R6835), .in2(6 'd 56));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op737 (.out1(_699), .in1(_698));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op738 (.out1(ck_idx_2605), .in1(R6834), .in2(_699));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2781 (.out1(R2782), .clock(clock), .in1(R2781));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2987 (.out1(R2988), .clock(clock), .in1(R2987));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3189 (.out1(R3190), .clock(clock), .in1(R3189));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3436 (.out1(R3437), .clock(clock), .in1(R3436));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3628 (.out1(R3629), .clock(clock), .in1(R3628));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3816 (.out1(R3817), .clock(clock), .in1(R3816));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4049 (.out1(R4050), .clock(clock), .in1(R4049));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4227 (.out1(R4228), .clock(clock), .in1(R4227));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4401 (.out1(R4402), .clock(clock), .in1(R4401));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4620 (.out1(R4621), .clock(clock), .in1(R4620));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4784 (.out1(R4785), .clock(clock), .in1(R4784));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4944 (.out1(R4945), .clock(clock), .in1(R4944));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5149 (.out1(R5150), .clock(clock), .in1(R5149));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5299 (.out1(R5300), .clock(clock), .in1(R5299));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5445 (.out1(R5446), .clock(clock), .in1(R5445));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5636 (.out1(R5637), .clock(clock), .in1(R5636));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5772 (.out1(R5773), .clock(clock), .in1(R5772));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5904 (.out1(R5905), .clock(clock), .in1(R5904));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6080 (.out1(R6081), .clock(clock), .in1(R6080));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6201 (.out1(R6202), .clock(clock), .in1(R6201));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6318 (.out1(R6319), .clock(clock), .in1(R6318));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6481 (.out1(R6482), .clock(clock), .in1(R6481));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6588 (.out1(R6589), .clock(clock), .in1(R6588));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6691 (.out1(R6692), .clock(clock), .in1(R6691));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6835 (.out1(R6836), .clock(clock), .in1(ck_idx_2605));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(4), .BITSIZE_out1(32), .PRECISION(32)) op739 (.out1(_700), .in1(R6836), .in2(4 'd 8));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op740 (.out1(_701), .in1(ip2_2595_D), .in2(6 'd 48));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2782 (.out1(R2783), .clock(clock), .in1(R2782));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2988 (.out1(R2989), .clock(clock), .in1(R2988));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3190 (.out1(R3191), .clock(clock), .in1(R3190));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3437 (.out1(R3438), .clock(clock), .in1(R3437));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3629 (.out1(R3630), .clock(clock), .in1(R3629));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3817 (.out1(R3818), .clock(clock), .in1(R3817));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4050 (.out1(R4051), .clock(clock), .in1(R4050));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4228 (.out1(R4229), .clock(clock), .in1(R4228));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4402 (.out1(R4403), .clock(clock), .in1(R4402));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4621 (.out1(R4622), .clock(clock), .in1(R4621));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4785 (.out1(R4786), .clock(clock), .in1(R4785));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4945 (.out1(R4946), .clock(clock), .in1(R4945));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5150 (.out1(R5151), .clock(clock), .in1(R5150));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5300 (.out1(R5301), .clock(clock), .in1(R5300));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5446 (.out1(R5447), .clock(clock), .in1(R5446));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5637 (.out1(R5638), .clock(clock), .in1(R5637));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5773 (.out1(R5774), .clock(clock), .in1(R5773));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5905 (.out1(R5906), .clock(clock), .in1(R5905));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6081 (.out1(R6082), .clock(clock), .in1(R6081));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6202 (.out1(R6203), .clock(clock), .in1(R6202));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6319 (.out1(R6320), .clock(clock), .in1(R6319));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6482 (.out1(R6483), .clock(clock), .in1(R6482));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6589 (.out1(R6590), .clock(clock), .in1(R6589));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6692 (.out1(R6693), .clock(clock), .in1(R6692));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6836 (.out1(R6837), .clock(clock), .in1(_700));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6837 (.out1(R6838), .clock(clock), .in1(_701));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op741 (.out1(_702), .in1(R6838));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(8), .BITSIZE_out1(32)) op742 (.out1(_703), .in1(_702), .in2(8 'd 255));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op743 (.out1(idx_sail_2606), .in1(R6837), .in2(_703));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(3), .BITSIZE_out1(32), .PRECISION(32)) op744 (.out1(idx_2607), .in1(idx_sail_2606), .in2(3 'd 6));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2783 (.out1(R2784), .clock(clock), .in1(R2783));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2989 (.out1(R2990), .clock(clock), .in1(R2989));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3191 (.out1(R3192), .clock(clock), .in1(R3191));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3438 (.out1(R3439), .clock(clock), .in1(R3438));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3630 (.out1(R3631), .clock(clock), .in1(R3630));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3818 (.out1(R3819), .clock(clock), .in1(R3818));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4051 (.out1(R4052), .clock(clock), .in1(R4051));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4229 (.out1(R4230), .clock(clock), .in1(R4229));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4403 (.out1(R4404), .clock(clock), .in1(R4403));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4622 (.out1(R4623), .clock(clock), .in1(R4622));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4786 (.out1(R4787), .clock(clock), .in1(R4786));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4946 (.out1(R4947), .clock(clock), .in1(R4946));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5151 (.out1(R5152), .clock(clock), .in1(R5151));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5301 (.out1(R5302), .clock(clock), .in1(R5301));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5447 (.out1(R5448), .clock(clock), .in1(R5447));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5638 (.out1(R5639), .clock(clock), .in1(R5638));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5774 (.out1(R5775), .clock(clock), .in1(R5774));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5906 (.out1(R5907), .clock(clock), .in1(R5906));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6082 (.out1(R6083), .clock(clock), .in1(R6082));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6203 (.out1(R6204), .clock(clock), .in1(R6203));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6320 (.out1(R6321), .clock(clock), .in1(R6320));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6483 (.out1(R6484), .clock(clock), .in1(R6483));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6590 (.out1(R6591), .clock(clock), .in1(R6590));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6693 (.out1(R6694), .clock(clock), .in1(R6693));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6838 (.out1(R6839), .clock(clock), .in1(idx_sail_2606));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6841 (.out1(R6842), .clock(clock), .in1(idx_2607));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op746 (.out1(_704), .in1(R6842));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op747 (.out1(_705), .in1(_704), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2784 (.out1(R2785), .clock(clock), .in1(R2784));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2990 (.out1(R2991), .clock(clock), .in1(R2990));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3192 (.out1(R3193), .clock(clock), .in1(R3192));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3439 (.out1(R3440), .clock(clock), .in1(R3439));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3631 (.out1(R3632), .clock(clock), .in1(R3631));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3819 (.out1(R3820), .clock(clock), .in1(R3819));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4052 (.out1(R4053), .clock(clock), .in1(R4052));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4230 (.out1(R4231), .clock(clock), .in1(R4230));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4404 (.out1(R4405), .clock(clock), .in1(R4404));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4623 (.out1(R4624), .clock(clock), .in1(R4623));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4787 (.out1(R4788), .clock(clock), .in1(R4787));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4947 (.out1(R4948), .clock(clock), .in1(R4947));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5152 (.out1(R5153), .clock(clock), .in1(R5152));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5302 (.out1(R5303), .clock(clock), .in1(R5302));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5448 (.out1(R5449), .clock(clock), .in1(R5448));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5639 (.out1(R5640), .clock(clock), .in1(R5639));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5775 (.out1(R5776), .clock(clock), .in1(R5775));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5907 (.out1(R5908), .clock(clock), .in1(R5907));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6083 (.out1(R6084), .clock(clock), .in1(R6083));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6204 (.out1(R6205), .clock(clock), .in1(R6204));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6321 (.out1(R6322), .clock(clock), .in1(R6321));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6484 (.out1(R6485), .clock(clock), .in1(R6484));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6591 (.out1(R6592), .clock(clock), .in1(R6591));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6694 (.out1(R6695), .clock(clock), .in1(R6694));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6839 (.out1(R6840), .clock(clock), .in1(R6839));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6842 (.out1(R6843), .clock(clock), .in1(R6842));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6934 (.out1(R6935), .clock(clock), .in1(_705));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op748 (.out1(_706), .in1(c80_bitmap_2609_D), .in2(R6935));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2785 (.out1(R2786), .clock(clock), .in1(R2785));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2991 (.out1(R2992), .clock(clock), .in1(R2991));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3193 (.out1(R3194), .clock(clock), .in1(R3193));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3440 (.out1(R3441), .clock(clock), .in1(R3440));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3632 (.out1(R3633), .clock(clock), .in1(R3632));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3820 (.out1(R3821), .clock(clock), .in1(R3820));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4053 (.out1(R4054), .clock(clock), .in1(R4053));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4231 (.out1(R4232), .clock(clock), .in1(R4231));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4405 (.out1(R4406), .clock(clock), .in1(R4405));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4624 (.out1(R4625), .clock(clock), .in1(R4624));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4788 (.out1(R4789), .clock(clock), .in1(R4788));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4948 (.out1(R4949), .clock(clock), .in1(R4948));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5153 (.out1(R5154), .clock(clock), .in1(R5153));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5303 (.out1(R5304), .clock(clock), .in1(R5303));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5449 (.out1(R5450), .clock(clock), .in1(R5449));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5640 (.out1(R5641), .clock(clock), .in1(R5640));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5776 (.out1(R5777), .clock(clock), .in1(R5776));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5908 (.out1(R5909), .clock(clock), .in1(R5908));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6084 (.out1(R6085), .clock(clock), .in1(R6084));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6205 (.out1(R6206), .clock(clock), .in1(R6205));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6322 (.out1(R6323), .clock(clock), .in1(R6322));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6485 (.out1(R6486), .clock(clock), .in1(R6485));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6592 (.out1(R6593), .clock(clock), .in1(R6592));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6695 (.out1(R6696), .clock(clock), .in1(R6695));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6840 (.out1(R6841), .clock(clock), .in1(R6840));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6843 (.out1(R6844), .clock(clock), .in1(R6843));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6935 (.out1(R6936), .clock(clock), .in1(_706));
  SRAM op749 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_707),.ADR(R6936));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op745 (.out1(off_2608), .in1(R6841), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op750 (.out1(_708), .in1(64 'd 9223372036854775808), .in2(off_2608));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2786 (.out1(R2787), .clock(clock), .in1(R2786));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2992 (.out1(R2993), .clock(clock), .in1(R2992));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3194 (.out1(R3195), .clock(clock), .in1(R3194));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3441 (.out1(R3442), .clock(clock), .in1(R3441));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3633 (.out1(R3634), .clock(clock), .in1(R3633));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3821 (.out1(R3822), .clock(clock), .in1(R3821));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4054 (.out1(R4055), .clock(clock), .in1(R4054));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4232 (.out1(R4233), .clock(clock), .in1(R4232));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4406 (.out1(R4407), .clock(clock), .in1(R4406));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4625 (.out1(R4626), .clock(clock), .in1(R4625));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4789 (.out1(R4790), .clock(clock), .in1(R4789));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4949 (.out1(R4950), .clock(clock), .in1(R4949));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5154 (.out1(R5155), .clock(clock), .in1(R5154));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5304 (.out1(R5305), .clock(clock), .in1(R5304));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5450 (.out1(R5451), .clock(clock), .in1(R5450));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5641 (.out1(R5642), .clock(clock), .in1(R5641));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5777 (.out1(R5778), .clock(clock), .in1(R5777));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5909 (.out1(R5910), .clock(clock), .in1(R5909));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6085 (.out1(R6086), .clock(clock), .in1(R6085));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6206 (.out1(R6207), .clock(clock), .in1(R6206));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6323 (.out1(R6324), .clock(clock), .in1(R6323));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6486 (.out1(R6487), .clock(clock), .in1(R6486));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6593 (.out1(R6594), .clock(clock), .in1(R6593));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6696 (.out1(R6697), .clock(clock), .in1(R6696));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6844 (.out1(R6845), .clock(clock), .in1(R6844));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6936 (.out1(R6937), .clock(clock), .in1(_707));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6937 (.out1(R6938), .clock(clock), .in1(off_2608));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7026 (.out1(R7027), .clock(clock), .in1(_708));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op751 (.out1(_709), .in1(R6937), .in2(R7027));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op752 (.out1(ifout752), .in1(_709), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op813 (.out1(_770), .in1(R6845));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op814 (.out1(_771), .in1(_770), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2787 (.out1(R2788), .clock(clock), .in1(R2787));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2993 (.out1(R2994), .clock(clock), .in1(R2993));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3195 (.out1(R3196), .clock(clock), .in1(R3195));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3442 (.out1(R3443), .clock(clock), .in1(R3442));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3634 (.out1(R3635), .clock(clock), .in1(R3634));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3822 (.out1(R3823), .clock(clock), .in1(R3822));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4055 (.out1(R4056), .clock(clock), .in1(R4055));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4233 (.out1(R4234), .clock(clock), .in1(R4233));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4407 (.out1(R4408), .clock(clock), .in1(R4407));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4626 (.out1(R4627), .clock(clock), .in1(R4626));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4790 (.out1(R4791), .clock(clock), .in1(R4790));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4950 (.out1(R4951), .clock(clock), .in1(R4950));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5155 (.out1(R5156), .clock(clock), .in1(R5155));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5305 (.out1(R5306), .clock(clock), .in1(R5305));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5451 (.out1(R5452), .clock(clock), .in1(R5451));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5642 (.out1(R5643), .clock(clock), .in1(R5642));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5778 (.out1(R5779), .clock(clock), .in1(R5778));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5910 (.out1(R5911), .clock(clock), .in1(R5910));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6086 (.out1(R6087), .clock(clock), .in1(R6086));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6207 (.out1(R6208), .clock(clock), .in1(R6207));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6324 (.out1(R6325), .clock(clock), .in1(R6324));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6487 (.out1(R6488), .clock(clock), .in1(R6487));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6594 (.out1(R6595), .clock(clock), .in1(R6594));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6697 (.out1(R6698), .clock(clock), .in1(R6697));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6845 (.out1(R6846), .clock(clock), .in1(R6845));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6938 (.out1(R6939), .clock(clock), .in1(R6938));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7027 (.out1(R7028), .clock(clock), .in1(ifout752));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7122 (.out1(R7123), .clock(clock), .in1(_771));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op807 (.out1(_764), .in1(R6846));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op797 (.out1(_754), .in1(R6846));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op791 (.out1(_748), .in1(R6846));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op779 (.out1(_736), .in1(R6846));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op773 (.out1(_730), .in1(R6846));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op763 (.out1(_720), .in1(R6846));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op808 (.out1(_765), .in1(_764), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op798 (.out1(_755), .in1(_754), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op792 (.out1(_749), .in1(_748), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op780 (.out1(_737), .in1(_736), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op774 (.out1(_731), .in1(_730), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op764 (.out1(_721), .in1(_720), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op815 (.out1(_772), .in1(c80_bitmap_2609_D), .in2(R7123));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2788 (.out1(R2789), .clock(clock), .in1(R2788));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2994 (.out1(R2995), .clock(clock), .in1(R2994));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3196 (.out1(R3197), .clock(clock), .in1(R3196));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3443 (.out1(R3444), .clock(clock), .in1(R3443));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3635 (.out1(R3636), .clock(clock), .in1(R3635));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3823 (.out1(R3824), .clock(clock), .in1(R3823));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4056 (.out1(R4057), .clock(clock), .in1(R4056));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4234 (.out1(R4235), .clock(clock), .in1(R4234));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4408 (.out1(R4409), .clock(clock), .in1(R4408));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4627 (.out1(R4628), .clock(clock), .in1(R4627));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4791 (.out1(R4792), .clock(clock), .in1(R4791));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4951 (.out1(R4952), .clock(clock), .in1(R4951));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5156 (.out1(R5157), .clock(clock), .in1(R5156));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5306 (.out1(R5307), .clock(clock), .in1(R5306));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5452 (.out1(R5453), .clock(clock), .in1(R5452));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5643 (.out1(R5644), .clock(clock), .in1(R5643));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5779 (.out1(R5780), .clock(clock), .in1(R5779));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5911 (.out1(R5912), .clock(clock), .in1(R5911));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6087 (.out1(R6088), .clock(clock), .in1(R6087));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6208 (.out1(R6209), .clock(clock), .in1(R6208));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6325 (.out1(R6326), .clock(clock), .in1(R6325));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6488 (.out1(R6489), .clock(clock), .in1(R6488));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6595 (.out1(R6596), .clock(clock), .in1(R6595));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6698 (.out1(R6699), .clock(clock), .in1(R6698));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6846 (.out1(R6847), .clock(clock), .in1(R6846));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6939 (.out1(R6940), .clock(clock), .in1(R6939));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7028 (.out1(R7029), .clock(clock), .in1(R7028));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7123 (.out1(R7124), .clock(clock), .in1(_765));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7124 (.out1(R7125), .clock(clock), .in1(_755));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7125 (.out1(R7126), .clock(clock), .in1(_749));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7126 (.out1(R7127), .clock(clock), .in1(_737));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7127 (.out1(R7128), .clock(clock), .in1(_731));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7128 (.out1(R7129), .clock(clock), .in1(_721));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7129 (.out1(R7130), .clock(clock), .in1(_772));
  SRAM op816 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_773),.ADR(R7130));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op757 (.out1(_714), .in1(R6847));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op758 (.out1(_715), .in1(_714), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op809 (.out1(_766), .in1(c80_bitmap_2609_D), .in2(R7124));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op799 (.out1(_756), .in1(c80_bitmap_2609_D), .in2(R7125));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op793 (.out1(_750), .in1(c80_bitmap_2609_D), .in2(R7126));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op781 (.out1(_738), .in1(c80_bitmap_2609_D), .in2(R7127));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op775 (.out1(_732), .in1(c80_bitmap_2609_D), .in2(R7128));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op765 (.out1(_722), .in1(c80_bitmap_2609_D), .in2(R7129));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2789 (.out1(R2790), .clock(clock), .in1(R2789));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2995 (.out1(R2996), .clock(clock), .in1(R2995));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3197 (.out1(R3198), .clock(clock), .in1(R3197));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3444 (.out1(R3445), .clock(clock), .in1(R3444));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3636 (.out1(R3637), .clock(clock), .in1(R3636));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3824 (.out1(R3825), .clock(clock), .in1(R3824));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4057 (.out1(R4058), .clock(clock), .in1(R4057));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4235 (.out1(R4236), .clock(clock), .in1(R4235));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4409 (.out1(R4410), .clock(clock), .in1(R4409));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4628 (.out1(R4629), .clock(clock), .in1(R4628));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4792 (.out1(R4793), .clock(clock), .in1(R4792));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4952 (.out1(R4953), .clock(clock), .in1(R4952));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5157 (.out1(R5158), .clock(clock), .in1(R5157));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5307 (.out1(R5308), .clock(clock), .in1(R5307));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5453 (.out1(R5454), .clock(clock), .in1(R5453));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5644 (.out1(R5645), .clock(clock), .in1(R5644));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5780 (.out1(R5781), .clock(clock), .in1(R5780));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5912 (.out1(R5913), .clock(clock), .in1(R5912));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6088 (.out1(R6089), .clock(clock), .in1(R6088));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6209 (.out1(R6210), .clock(clock), .in1(R6209));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6326 (.out1(R6327), .clock(clock), .in1(R6326));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6489 (.out1(R6490), .clock(clock), .in1(R6489));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6596 (.out1(R6597), .clock(clock), .in1(R6596));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6699 (.out1(R6700), .clock(clock), .in1(R6699));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6847 (.out1(R6848), .clock(clock), .in1(R6847));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6940 (.out1(R6941), .clock(clock), .in1(R6940));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7029 (.out1(R7030), .clock(clock), .in1(R7029));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7130 (.out1(R7131), .clock(clock), .in1(_773));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7131 (.out1(R7132), .clock(clock), .in1(_715));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7132 (.out1(R7133), .clock(clock), .in1(_766));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7133 (.out1(R7134), .clock(clock), .in1(_756));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7134 (.out1(R7135), .clock(clock), .in1(_750));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7135 (.out1(R7136), .clock(clock), .in1(_738));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7136 (.out1(R7137), .clock(clock), .in1(_732));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7137 (.out1(R7138), .clock(clock), .in1(_722));
  SRAM op810 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_767),.ADR(R7133));
  SRAM op800 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_757),.ADR(R7134));
  SRAM op794 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_751),.ADR(R7135));
  SRAM op782 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_739),.ADR(R7136));
  SRAM op776 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_733),.ADR(R7137));
  SRAM op766 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_723),.ADR(R7138));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op817 (.out1(_774), .in1(7 'd 64), .in2(R6941));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op759 (.out1(_716), .in1(c80_bitmap_2609_D), .in2(R7132));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op818 (.out1(_775), .in1(R7131), .in2(_774));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op811 (.out1(_768), .in1(7 'd 64), .in2(R6941));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op801 (.out1(_758), .in1(7 'd 64), .in2(R6941));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op783 (.out1(_740), .in1(7 'd 64), .in2(R6941));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2790 (.out1(R2791), .clock(clock), .in1(R2790));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2996 (.out1(R2997), .clock(clock), .in1(R2996));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3198 (.out1(R3199), .clock(clock), .in1(R3198));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3445 (.out1(R3446), .clock(clock), .in1(R3445));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3637 (.out1(R3638), .clock(clock), .in1(R3637));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3825 (.out1(R3826), .clock(clock), .in1(R3825));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4058 (.out1(R4059), .clock(clock), .in1(R4058));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4236 (.out1(R4237), .clock(clock), .in1(R4236));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4410 (.out1(R4411), .clock(clock), .in1(R4410));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4629 (.out1(R4630), .clock(clock), .in1(R4629));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4793 (.out1(R4794), .clock(clock), .in1(R4793));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4953 (.out1(R4954), .clock(clock), .in1(R4953));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5158 (.out1(R5159), .clock(clock), .in1(R5158));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5308 (.out1(R5309), .clock(clock), .in1(R5308));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5454 (.out1(R5455), .clock(clock), .in1(R5454));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5645 (.out1(R5646), .clock(clock), .in1(R5645));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5781 (.out1(R5782), .clock(clock), .in1(R5781));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5913 (.out1(R5914), .clock(clock), .in1(R5913));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6089 (.out1(R6090), .clock(clock), .in1(R6089));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6210 (.out1(R6211), .clock(clock), .in1(R6210));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6327 (.out1(R6328), .clock(clock), .in1(R6327));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6490 (.out1(R6491), .clock(clock), .in1(R6490));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6597 (.out1(R6598), .clock(clock), .in1(R6597));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6700 (.out1(R6701), .clock(clock), .in1(R6700));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6848 (.out1(R6849), .clock(clock), .in1(R6848));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6941 (.out1(R6942), .clock(clock), .in1(R6941));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7030 (.out1(R7031), .clock(clock), .in1(R7030));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7138 (.out1(R7139), .clock(clock), .in1(_767));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7139 (.out1(R7140), .clock(clock), .in1(_757));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7140 (.out1(R7141), .clock(clock), .in1(_751));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7141 (.out1(R7142), .clock(clock), .in1(_739));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7142 (.out1(R7143), .clock(clock), .in1(_733));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7143 (.out1(R7144), .clock(clock), .in1(_723));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7144 (.out1(R7145), .clock(clock), .in1(_716));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7145 (.out1(R7146), .clock(clock), .in1(_775));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7146 (.out1(R7147), .clock(clock), .in1(_768));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7147 (.out1(R7148), .clock(clock), .in1(_758));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7148 (.out1(R7149), .clock(clock), .in1(_740));
  SRAM op760 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_717),.ADR(R7145));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op819 (.out1(_776), .in1(R7146), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op812 (.out1(_769), .in1(R7139), .in2(R7147));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op802 (.out1(_759), .in1(R7140), .in2(R7148));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op795 (.out1(_752), .in1(7 'd 64), .in2(R6942));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op784 (.out1(_741), .in1(R7142), .in2(R7149));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op777 (.out1(_734), .in1(7 'd 64), .in2(R6942));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op767 (.out1(_724), .in1(7 'd 64), .in2(R6942));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op820 (.out1(_777), .in1(_776), .in2(63 'd 6148914691236517205));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op821 (.out1(_778), .in1(_769), .in2(_777));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op803 (.out1(_760), .in1(_759), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op796 (.out1(_753), .in1(R7141), .in2(_752));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op785 (.out1(_742), .in1(_741), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op778 (.out1(_735), .in1(R7143), .in2(_734));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op768 (.out1(_725), .in1(R7144), .in2(_724));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op761 (.out1(_718), .in1(7 'd 64), .in2(R6942));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2791 (.out1(R2792), .clock(clock), .in1(R2791));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2997 (.out1(R2998), .clock(clock), .in1(R2997));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3199 (.out1(R3200), .clock(clock), .in1(R3199));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3446 (.out1(R3447), .clock(clock), .in1(R3446));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3638 (.out1(R3639), .clock(clock), .in1(R3638));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3826 (.out1(R3827), .clock(clock), .in1(R3826));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4059 (.out1(R4060), .clock(clock), .in1(R4059));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4237 (.out1(R4238), .clock(clock), .in1(R4237));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4411 (.out1(R4412), .clock(clock), .in1(R4411));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4630 (.out1(R4631), .clock(clock), .in1(R4630));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4794 (.out1(R4795), .clock(clock), .in1(R4794));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4954 (.out1(R4955), .clock(clock), .in1(R4954));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5159 (.out1(R5160), .clock(clock), .in1(R5159));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5309 (.out1(R5310), .clock(clock), .in1(R5309));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5455 (.out1(R5456), .clock(clock), .in1(R5455));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5646 (.out1(R5647), .clock(clock), .in1(R5646));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5782 (.out1(R5783), .clock(clock), .in1(R5782));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5914 (.out1(R5915), .clock(clock), .in1(R5914));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6090 (.out1(R6091), .clock(clock), .in1(R6090));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6211 (.out1(R6212), .clock(clock), .in1(R6211));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6328 (.out1(R6329), .clock(clock), .in1(R6328));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6491 (.out1(R6492), .clock(clock), .in1(R6491));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6598 (.out1(R6599), .clock(clock), .in1(R6598));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6701 (.out1(R6702), .clock(clock), .in1(R6701));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6849 (.out1(R6850), .clock(clock), .in1(R6849));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6942 (.out1(R6943), .clock(clock), .in1(R6942));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7031 (.out1(R7032), .clock(clock), .in1(R7031));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7149 (.out1(R7150), .clock(clock), .in1(_717));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7150 (.out1(R7151), .clock(clock), .in1(_778));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7151 (.out1(R7152), .clock(clock), .in1(_760));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7152 (.out1(R7153), .clock(clock), .in1(_753));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7153 (.out1(R7154), .clock(clock), .in1(_742));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7154 (.out1(R7155), .clock(clock), .in1(_735));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7155 (.out1(R7156), .clock(clock), .in1(_725));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7156 (.out1(R7157), .clock(clock), .in1(_718));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op753 (.out1(_710), .in1(R6850));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op804 (.out1(_761), .in1(R7152), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op822 (.out1(_779), .in1(R7151), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op805 (.out1(_762), .in1(R7153), .in2(_761));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op786 (.out1(_743), .in1(R7154), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op769 (.out1(_726), .in1(R7156), .in2(1 'd 1));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op787 (.out1(_744), .in1(R7155), .in2(_743));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op762 (.out1(_719), .in1(R7150), .in2(R7157));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op754 (.out1(_711), .in1(_710), .in2(2 'd 2));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op823 (.out1(_780), .in1(_779), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op806 (.out1(_763), .in1(_762), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op770 (.out1(_727), .in1(_726), .in2(63 'd 6148914691236517205));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op824 (.out1(_781), .in1(_763), .in2(_780));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op788 (.out1(_745), .in1(_744), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op771 (.out1(_728), .in1(_719), .in2(_727));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2792 (.out1(R2793), .clock(clock), .in1(R2792));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2998 (.out1(R2999), .clock(clock), .in1(R2998));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3200 (.out1(R3201), .clock(clock), .in1(R3200));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3447 (.out1(R3448), .clock(clock), .in1(R3447));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3639 (.out1(R3640), .clock(clock), .in1(R3639));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3827 (.out1(R3828), .clock(clock), .in1(R3827));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4060 (.out1(R4061), .clock(clock), .in1(R4060));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4238 (.out1(R4239), .clock(clock), .in1(R4238));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4412 (.out1(R4413), .clock(clock), .in1(R4412));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4631 (.out1(R4632), .clock(clock), .in1(R4631));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4795 (.out1(R4796), .clock(clock), .in1(R4795));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4955 (.out1(R4956), .clock(clock), .in1(R4955));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5160 (.out1(R5161), .clock(clock), .in1(R5160));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5310 (.out1(R5311), .clock(clock), .in1(R5310));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5456 (.out1(R5457), .clock(clock), .in1(R5456));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5647 (.out1(R5648), .clock(clock), .in1(R5647));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5783 (.out1(R5784), .clock(clock), .in1(R5783));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5915 (.out1(R5916), .clock(clock), .in1(R5915));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6091 (.out1(R6092), .clock(clock), .in1(R6091));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6212 (.out1(R6213), .clock(clock), .in1(R6212));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6329 (.out1(R6330), .clock(clock), .in1(R6329));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6492 (.out1(R6493), .clock(clock), .in1(R6492));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6599 (.out1(R6600), .clock(clock), .in1(R6599));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6702 (.out1(R6703), .clock(clock), .in1(R6702));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6850 (.out1(R6851), .clock(clock), .in1(R6850));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6943 (.out1(R6944), .clock(clock), .in1(R6943));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7032 (.out1(R7033), .clock(clock), .in1(R7032));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7157 (.out1(R7158), .clock(clock), .in1(_711));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7158 (.out1(R7159), .clock(clock), .in1(_781));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7159 (.out1(R7160), .clock(clock), .in1(_745));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7160 (.out1(R7161), .clock(clock), .in1(_728));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op789 (.out1(_746), .in1(R7160), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op772 (.out1(_729), .in1(R7161), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op825 (.out1(_782), .in1(R7159), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op790 (.out1(_747), .in1(_729), .in2(_746));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op755 (.out1(_712), .in1(c80_popcnt_2614_D), .in2(R7158));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op826 (.out1(_783), .in1(_747), .in2(_782));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op827 (.out1(_784), .in1(_783), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2793 (.out1(R2794), .clock(clock), .in1(R2793));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2999 (.out1(R3000), .clock(clock), .in1(R2999));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3201 (.out1(R3202), .clock(clock), .in1(R3201));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3448 (.out1(R3449), .clock(clock), .in1(R3448));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3640 (.out1(R3641), .clock(clock), .in1(R3640));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3828 (.out1(R3829), .clock(clock), .in1(R3828));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4061 (.out1(R4062), .clock(clock), .in1(R4061));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4239 (.out1(R4240), .clock(clock), .in1(R4239));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4413 (.out1(R4414), .clock(clock), .in1(R4413));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4632 (.out1(R4633), .clock(clock), .in1(R4632));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4796 (.out1(R4797), .clock(clock), .in1(R4796));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4956 (.out1(R4957), .clock(clock), .in1(R4956));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5161 (.out1(R5162), .clock(clock), .in1(R5161));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5311 (.out1(R5312), .clock(clock), .in1(R5311));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5457 (.out1(R5458), .clock(clock), .in1(R5457));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5648 (.out1(R5649), .clock(clock), .in1(R5648));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5784 (.out1(R5785), .clock(clock), .in1(R5784));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5916 (.out1(R5917), .clock(clock), .in1(R5916));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6092 (.out1(R6093), .clock(clock), .in1(R6092));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6213 (.out1(R6214), .clock(clock), .in1(R6213));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6330 (.out1(R6331), .clock(clock), .in1(R6330));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6493 (.out1(R6494), .clock(clock), .in1(R6493));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6600 (.out1(R6601), .clock(clock), .in1(R6600));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6703 (.out1(R6704), .clock(clock), .in1(R6703));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6851 (.out1(R6852), .clock(clock), .in1(R6851));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6944 (.out1(R6945), .clock(clock), .in1(R6944));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7033 (.out1(R7034), .clock(clock), .in1(R7033));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7161 (.out1(R7162), .clock(clock), .in1(_712));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7162 (.out1(R7163), .clock(clock), .in1(_784));
  SRAM op756 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_713),.ADR(R7162));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op828 (.out1(_785), .in1(R7163), .in2(57 'd 72340172838076673));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2794 (.out1(R2795), .clock(clock), .in1(R2794));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3000 (.out1(R3001), .clock(clock), .in1(R3000));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3202 (.out1(R3203), .clock(clock), .in1(R3202));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3449 (.out1(R3450), .clock(clock), .in1(R3449));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3641 (.out1(R3642), .clock(clock), .in1(R3641));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3829 (.out1(R3830), .clock(clock), .in1(R3829));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4062 (.out1(R4063), .clock(clock), .in1(R4062));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4240 (.out1(R4241), .clock(clock), .in1(R4240));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4414 (.out1(R4415), .clock(clock), .in1(R4414));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4633 (.out1(R4634), .clock(clock), .in1(R4633));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4797 (.out1(R4798), .clock(clock), .in1(R4797));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4957 (.out1(R4958), .clock(clock), .in1(R4957));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5162 (.out1(R5163), .clock(clock), .in1(R5162));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5312 (.out1(R5313), .clock(clock), .in1(R5312));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5458 (.out1(R5459), .clock(clock), .in1(R5458));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5649 (.out1(R5650), .clock(clock), .in1(R5649));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5785 (.out1(R5786), .clock(clock), .in1(R5785));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5917 (.out1(R5918), .clock(clock), .in1(R5917));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6093 (.out1(R6094), .clock(clock), .in1(R6093));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6214 (.out1(R6215), .clock(clock), .in1(R6214));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6331 (.out1(R6332), .clock(clock), .in1(R6331));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6494 (.out1(R6495), .clock(clock), .in1(R6494));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6601 (.out1(R6602), .clock(clock), .in1(R6601));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6704 (.out1(R6705), .clock(clock), .in1(R6704));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6852 (.out1(R6853), .clock(clock), .in1(R6852));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6945 (.out1(R6946), .clock(clock), .in1(R6945));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7034 (.out1(R7035), .clock(clock), .in1(R7034));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7163 (.out1(R7164), .clock(clock), .in1(_713));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7164 (.out1(R7165), .clock(clock), .in1(_785));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op829 (.out1(_786), .in1(R7165), .in2(6 'd 56));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op830 (.out1(_787), .in1(_786));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op831 (.out1(ck_idx_2615), .in1(R7164), .in2(_787));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2795 (.out1(R2796), .clock(clock), .in1(R2795));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3001 (.out1(R3002), .clock(clock), .in1(R3001));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3203 (.out1(R3204), .clock(clock), .in1(R3203));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3450 (.out1(R3451), .clock(clock), .in1(R3450));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3642 (.out1(R3643), .clock(clock), .in1(R3642));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3830 (.out1(R3831), .clock(clock), .in1(R3830));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4063 (.out1(R4064), .clock(clock), .in1(R4063));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4241 (.out1(R4242), .clock(clock), .in1(R4241));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4415 (.out1(R4416), .clock(clock), .in1(R4415));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4634 (.out1(R4635), .clock(clock), .in1(R4634));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4798 (.out1(R4799), .clock(clock), .in1(R4798));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4958 (.out1(R4959), .clock(clock), .in1(R4958));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5163 (.out1(R5164), .clock(clock), .in1(R5163));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5313 (.out1(R5314), .clock(clock), .in1(R5313));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5459 (.out1(R5460), .clock(clock), .in1(R5459));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5650 (.out1(R5651), .clock(clock), .in1(R5650));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5786 (.out1(R5787), .clock(clock), .in1(R5786));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5918 (.out1(R5919), .clock(clock), .in1(R5918));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6094 (.out1(R6095), .clock(clock), .in1(R6094));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6215 (.out1(R6216), .clock(clock), .in1(R6215));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6332 (.out1(R6333), .clock(clock), .in1(R6332));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6495 (.out1(R6496), .clock(clock), .in1(R6495));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6602 (.out1(R6603), .clock(clock), .in1(R6602));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6705 (.out1(R6706), .clock(clock), .in1(R6705));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6853 (.out1(R6854), .clock(clock), .in1(R6853));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6946 (.out1(R6947), .clock(clock), .in1(R6946));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7035 (.out1(R7036), .clock(clock), .in1(R7035));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7165 (.out1(R7166), .clock(clock), .in1(ck_idx_2615));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(4), .BITSIZE_out1(32), .PRECISION(32)) op832 (.out1(_788), .in1(R7166), .in2(4 'd 8));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op833 (.out1(_789), .in1(ip2_2595_D), .in2(6 'd 40));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2796 (.out1(R2797), .clock(clock), .in1(R2796));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3002 (.out1(R3003), .clock(clock), .in1(R3002));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3204 (.out1(R3205), .clock(clock), .in1(R3204));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3451 (.out1(R3452), .clock(clock), .in1(R3451));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3643 (.out1(R3644), .clock(clock), .in1(R3643));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3831 (.out1(R3832), .clock(clock), .in1(R3831));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4064 (.out1(R4065), .clock(clock), .in1(R4064));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4242 (.out1(R4243), .clock(clock), .in1(R4242));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4416 (.out1(R4417), .clock(clock), .in1(R4416));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4635 (.out1(R4636), .clock(clock), .in1(R4635));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4799 (.out1(R4800), .clock(clock), .in1(R4799));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4959 (.out1(R4960), .clock(clock), .in1(R4959));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5164 (.out1(R5165), .clock(clock), .in1(R5164));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5314 (.out1(R5315), .clock(clock), .in1(R5314));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5460 (.out1(R5461), .clock(clock), .in1(R5460));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5651 (.out1(R5652), .clock(clock), .in1(R5651));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5787 (.out1(R5788), .clock(clock), .in1(R5787));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5919 (.out1(R5920), .clock(clock), .in1(R5919));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6095 (.out1(R6096), .clock(clock), .in1(R6095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6216 (.out1(R6217), .clock(clock), .in1(R6216));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6333 (.out1(R6334), .clock(clock), .in1(R6333));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6496 (.out1(R6497), .clock(clock), .in1(R6496));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6603 (.out1(R6604), .clock(clock), .in1(R6603));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6706 (.out1(R6707), .clock(clock), .in1(R6706));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6854 (.out1(R6855), .clock(clock), .in1(R6854));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6947 (.out1(R6948), .clock(clock), .in1(R6947));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7036 (.out1(R7037), .clock(clock), .in1(R7036));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7166 (.out1(R7167), .clock(clock), .in1(_788));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7167 (.out1(R7168), .clock(clock), .in1(_789));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op834 (.out1(_790), .in1(R7168));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(8), .BITSIZE_out1(32)) op835 (.out1(_791), .in1(_790), .in2(8 'd 255));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op836 (.out1(idx_sail_2616), .in1(R7167), .in2(_791));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(3), .BITSIZE_out1(32), .PRECISION(32)) op837 (.out1(idx_2617), .in1(idx_sail_2616), .in2(3 'd 6));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2797 (.out1(R2798), .clock(clock), .in1(R2797));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3003 (.out1(R3004), .clock(clock), .in1(R3003));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3205 (.out1(R3206), .clock(clock), .in1(R3205));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3452 (.out1(R3453), .clock(clock), .in1(R3452));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3644 (.out1(R3645), .clock(clock), .in1(R3644));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3832 (.out1(R3833), .clock(clock), .in1(R3832));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4065 (.out1(R4066), .clock(clock), .in1(R4065));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4243 (.out1(R4244), .clock(clock), .in1(R4243));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4417 (.out1(R4418), .clock(clock), .in1(R4417));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4636 (.out1(R4637), .clock(clock), .in1(R4636));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4800 (.out1(R4801), .clock(clock), .in1(R4800));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4960 (.out1(R4961), .clock(clock), .in1(R4960));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5165 (.out1(R5166), .clock(clock), .in1(R5165));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5315 (.out1(R5316), .clock(clock), .in1(R5315));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5461 (.out1(R5462), .clock(clock), .in1(R5461));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5652 (.out1(R5653), .clock(clock), .in1(R5652));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5788 (.out1(R5789), .clock(clock), .in1(R5788));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5920 (.out1(R5921), .clock(clock), .in1(R5920));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6096 (.out1(R6097), .clock(clock), .in1(R6096));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6217 (.out1(R6218), .clock(clock), .in1(R6217));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6334 (.out1(R6335), .clock(clock), .in1(R6334));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6497 (.out1(R6498), .clock(clock), .in1(R6497));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6604 (.out1(R6605), .clock(clock), .in1(R6604));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6707 (.out1(R6708), .clock(clock), .in1(R6707));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6855 (.out1(R6856), .clock(clock), .in1(R6855));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6948 (.out1(R6949), .clock(clock), .in1(R6948));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7037 (.out1(R7038), .clock(clock), .in1(R7037));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7168 (.out1(R7169), .clock(clock), .in1(idx_sail_2616));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7171 (.out1(R7172), .clock(clock), .in1(idx_2617));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op839 (.out1(_792), .in1(R7172));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op840 (.out1(_793), .in1(_792), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2798 (.out1(R2799), .clock(clock), .in1(R2798));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3004 (.out1(R3005), .clock(clock), .in1(R3004));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3206 (.out1(R3207), .clock(clock), .in1(R3206));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3453 (.out1(R3454), .clock(clock), .in1(R3453));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3645 (.out1(R3646), .clock(clock), .in1(R3645));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3833 (.out1(R3834), .clock(clock), .in1(R3833));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4066 (.out1(R4067), .clock(clock), .in1(R4066));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4244 (.out1(R4245), .clock(clock), .in1(R4244));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4418 (.out1(R4419), .clock(clock), .in1(R4418));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4637 (.out1(R4638), .clock(clock), .in1(R4637));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4801 (.out1(R4802), .clock(clock), .in1(R4801));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4961 (.out1(R4962), .clock(clock), .in1(R4961));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5166 (.out1(R5167), .clock(clock), .in1(R5166));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5316 (.out1(R5317), .clock(clock), .in1(R5316));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5462 (.out1(R5463), .clock(clock), .in1(R5462));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5653 (.out1(R5654), .clock(clock), .in1(R5653));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5789 (.out1(R5790), .clock(clock), .in1(R5789));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5921 (.out1(R5922), .clock(clock), .in1(R5921));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6097 (.out1(R6098), .clock(clock), .in1(R6097));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6218 (.out1(R6219), .clock(clock), .in1(R6218));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6335 (.out1(R6336), .clock(clock), .in1(R6335));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6498 (.out1(R6499), .clock(clock), .in1(R6498));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6605 (.out1(R6606), .clock(clock), .in1(R6605));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6708 (.out1(R6709), .clock(clock), .in1(R6708));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6856 (.out1(R6857), .clock(clock), .in1(R6856));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6949 (.out1(R6950), .clock(clock), .in1(R6949));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7038 (.out1(R7039), .clock(clock), .in1(R7038));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7169 (.out1(R7170), .clock(clock), .in1(R7169));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7172 (.out1(R7173), .clock(clock), .in1(R7172));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7250 (.out1(R7251), .clock(clock), .in1(_793));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op841 (.out1(_794), .in1(c88_bitmap_2619_D), .in2(R7251));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2799 (.out1(R2800), .clock(clock), .in1(R2799));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3005 (.out1(R3006), .clock(clock), .in1(R3005));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3207 (.out1(R3208), .clock(clock), .in1(R3207));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3454 (.out1(R3455), .clock(clock), .in1(R3454));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3646 (.out1(R3647), .clock(clock), .in1(R3646));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3834 (.out1(R3835), .clock(clock), .in1(R3834));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4067 (.out1(R4068), .clock(clock), .in1(R4067));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4245 (.out1(R4246), .clock(clock), .in1(R4245));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4419 (.out1(R4420), .clock(clock), .in1(R4419));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4638 (.out1(R4639), .clock(clock), .in1(R4638));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4802 (.out1(R4803), .clock(clock), .in1(R4802));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4962 (.out1(R4963), .clock(clock), .in1(R4962));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5167 (.out1(R5168), .clock(clock), .in1(R5167));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5317 (.out1(R5318), .clock(clock), .in1(R5317));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5463 (.out1(R5464), .clock(clock), .in1(R5463));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5654 (.out1(R5655), .clock(clock), .in1(R5654));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5790 (.out1(R5791), .clock(clock), .in1(R5790));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5922 (.out1(R5923), .clock(clock), .in1(R5922));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6098 (.out1(R6099), .clock(clock), .in1(R6098));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6219 (.out1(R6220), .clock(clock), .in1(R6219));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6336 (.out1(R6337), .clock(clock), .in1(R6336));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6499 (.out1(R6500), .clock(clock), .in1(R6499));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6606 (.out1(R6607), .clock(clock), .in1(R6606));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6709 (.out1(R6710), .clock(clock), .in1(R6709));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6857 (.out1(R6858), .clock(clock), .in1(R6857));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6950 (.out1(R6951), .clock(clock), .in1(R6950));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7039 (.out1(R7040), .clock(clock), .in1(R7039));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7170 (.out1(R7171), .clock(clock), .in1(R7170));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7173 (.out1(R7174), .clock(clock), .in1(R7173));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7251 (.out1(R7252), .clock(clock), .in1(_794));
  SRAM op842 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_795),.ADR(R7252));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op838 (.out1(off_2618), .in1(R7171), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op843 (.out1(_796), .in1(64 'd 9223372036854775808), .in2(off_2618));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2800 (.out1(R2801), .clock(clock), .in1(R2800));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3006 (.out1(R3007), .clock(clock), .in1(R3006));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3208 (.out1(R3209), .clock(clock), .in1(R3208));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3455 (.out1(R3456), .clock(clock), .in1(R3455));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3647 (.out1(R3648), .clock(clock), .in1(R3647));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3835 (.out1(R3836), .clock(clock), .in1(R3835));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4068 (.out1(R4069), .clock(clock), .in1(R4068));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4246 (.out1(R4247), .clock(clock), .in1(R4246));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4420 (.out1(R4421), .clock(clock), .in1(R4420));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4639 (.out1(R4640), .clock(clock), .in1(R4639));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4803 (.out1(R4804), .clock(clock), .in1(R4803));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4963 (.out1(R4964), .clock(clock), .in1(R4963));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5168 (.out1(R5169), .clock(clock), .in1(R5168));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5318 (.out1(R5319), .clock(clock), .in1(R5318));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5464 (.out1(R5465), .clock(clock), .in1(R5464));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5655 (.out1(R5656), .clock(clock), .in1(R5655));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5791 (.out1(R5792), .clock(clock), .in1(R5791));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5923 (.out1(R5924), .clock(clock), .in1(R5923));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6099 (.out1(R6100), .clock(clock), .in1(R6099));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6220 (.out1(R6221), .clock(clock), .in1(R6220));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6337 (.out1(R6338), .clock(clock), .in1(R6337));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6500 (.out1(R6501), .clock(clock), .in1(R6500));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6607 (.out1(R6608), .clock(clock), .in1(R6607));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6710 (.out1(R6711), .clock(clock), .in1(R6710));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6858 (.out1(R6859), .clock(clock), .in1(R6858));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6951 (.out1(R6952), .clock(clock), .in1(R6951));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7040 (.out1(R7041), .clock(clock), .in1(R7040));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7174 (.out1(R7175), .clock(clock), .in1(R7174));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7252 (.out1(R7253), .clock(clock), .in1(_795));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7253 (.out1(R7254), .clock(clock), .in1(off_2618));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7328 (.out1(R7329), .clock(clock), .in1(_796));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op844 (.out1(_797), .in1(R7253), .in2(R7329));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op845 (.out1(ifout845), .in1(_797), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op906 (.out1(_858), .in1(R7175));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op907 (.out1(_859), .in1(_858), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2801 (.out1(R2802), .clock(clock), .in1(R2801));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3007 (.out1(R3008), .clock(clock), .in1(R3007));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3209 (.out1(R3210), .clock(clock), .in1(R3209));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3456 (.out1(R3457), .clock(clock), .in1(R3456));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3648 (.out1(R3649), .clock(clock), .in1(R3648));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3836 (.out1(R3837), .clock(clock), .in1(R3836));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4069 (.out1(R4070), .clock(clock), .in1(R4069));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4247 (.out1(R4248), .clock(clock), .in1(R4247));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4421 (.out1(R4422), .clock(clock), .in1(R4421));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4640 (.out1(R4641), .clock(clock), .in1(R4640));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4804 (.out1(R4805), .clock(clock), .in1(R4804));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4964 (.out1(R4965), .clock(clock), .in1(R4964));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5169 (.out1(R5170), .clock(clock), .in1(R5169));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5319 (.out1(R5320), .clock(clock), .in1(R5319));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5465 (.out1(R5466), .clock(clock), .in1(R5465));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5656 (.out1(R5657), .clock(clock), .in1(R5656));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5792 (.out1(R5793), .clock(clock), .in1(R5792));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5924 (.out1(R5925), .clock(clock), .in1(R5924));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6100 (.out1(R6101), .clock(clock), .in1(R6100));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6221 (.out1(R6222), .clock(clock), .in1(R6221));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6338 (.out1(R6339), .clock(clock), .in1(R6338));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6501 (.out1(R6502), .clock(clock), .in1(R6501));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6608 (.out1(R6609), .clock(clock), .in1(R6608));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6711 (.out1(R6712), .clock(clock), .in1(R6711));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6859 (.out1(R6860), .clock(clock), .in1(R6859));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6952 (.out1(R6953), .clock(clock), .in1(R6952));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7041 (.out1(R7042), .clock(clock), .in1(R7041));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7175 (.out1(R7176), .clock(clock), .in1(R7175));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7254 (.out1(R7255), .clock(clock), .in1(R7254));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7329 (.out1(R7330), .clock(clock), .in1(ifout845));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7410 (.out1(R7411), .clock(clock), .in1(_859));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op900 (.out1(_852), .in1(R7176));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op890 (.out1(_842), .in1(R7176));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op884 (.out1(_836), .in1(R7176));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op872 (.out1(_824), .in1(R7176));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op866 (.out1(_818), .in1(R7176));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op856 (.out1(_808), .in1(R7176));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op901 (.out1(_853), .in1(_852), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op891 (.out1(_843), .in1(_842), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op885 (.out1(_837), .in1(_836), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op873 (.out1(_825), .in1(_824), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op867 (.out1(_819), .in1(_818), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op857 (.out1(_809), .in1(_808), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op908 (.out1(_860), .in1(c88_bitmap_2619_D), .in2(R7411));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2802 (.out1(R2803), .clock(clock), .in1(R2802));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3008 (.out1(R3009), .clock(clock), .in1(R3008));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3210 (.out1(R3211), .clock(clock), .in1(R3210));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3457 (.out1(R3458), .clock(clock), .in1(R3457));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3649 (.out1(R3650), .clock(clock), .in1(R3649));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3837 (.out1(R3838), .clock(clock), .in1(R3837));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4070 (.out1(R4071), .clock(clock), .in1(R4070));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4248 (.out1(R4249), .clock(clock), .in1(R4248));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4422 (.out1(R4423), .clock(clock), .in1(R4422));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4641 (.out1(R4642), .clock(clock), .in1(R4641));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4805 (.out1(R4806), .clock(clock), .in1(R4805));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4965 (.out1(R4966), .clock(clock), .in1(R4965));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5170 (.out1(R5171), .clock(clock), .in1(R5170));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5320 (.out1(R5321), .clock(clock), .in1(R5320));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5466 (.out1(R5467), .clock(clock), .in1(R5466));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5657 (.out1(R5658), .clock(clock), .in1(R5657));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5793 (.out1(R5794), .clock(clock), .in1(R5793));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5925 (.out1(R5926), .clock(clock), .in1(R5925));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6101 (.out1(R6102), .clock(clock), .in1(R6101));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6222 (.out1(R6223), .clock(clock), .in1(R6222));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6339 (.out1(R6340), .clock(clock), .in1(R6339));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6502 (.out1(R6503), .clock(clock), .in1(R6502));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6609 (.out1(R6610), .clock(clock), .in1(R6609));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6712 (.out1(R6713), .clock(clock), .in1(R6712));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6860 (.out1(R6861), .clock(clock), .in1(R6860));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6953 (.out1(R6954), .clock(clock), .in1(R6953));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7042 (.out1(R7043), .clock(clock), .in1(R7042));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7176 (.out1(R7177), .clock(clock), .in1(R7176));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7255 (.out1(R7256), .clock(clock), .in1(R7255));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7330 (.out1(R7331), .clock(clock), .in1(R7330));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7411 (.out1(R7412), .clock(clock), .in1(_853));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7412 (.out1(R7413), .clock(clock), .in1(_843));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7413 (.out1(R7414), .clock(clock), .in1(_837));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7414 (.out1(R7415), .clock(clock), .in1(_825));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7415 (.out1(R7416), .clock(clock), .in1(_819));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7416 (.out1(R7417), .clock(clock), .in1(_809));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7417 (.out1(R7418), .clock(clock), .in1(_860));
  SRAM op909 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_861),.ADR(R7418));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op850 (.out1(_802), .in1(R7177));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op851 (.out1(_803), .in1(_802), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op902 (.out1(_854), .in1(c88_bitmap_2619_D), .in2(R7412));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op892 (.out1(_844), .in1(c88_bitmap_2619_D), .in2(R7413));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op886 (.out1(_838), .in1(c88_bitmap_2619_D), .in2(R7414));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op874 (.out1(_826), .in1(c88_bitmap_2619_D), .in2(R7415));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op868 (.out1(_820), .in1(c88_bitmap_2619_D), .in2(R7416));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op858 (.out1(_810), .in1(c88_bitmap_2619_D), .in2(R7417));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2803 (.out1(R2804), .clock(clock), .in1(R2803));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3009 (.out1(R3010), .clock(clock), .in1(R3009));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3211 (.out1(R3212), .clock(clock), .in1(R3211));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3458 (.out1(R3459), .clock(clock), .in1(R3458));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3650 (.out1(R3651), .clock(clock), .in1(R3650));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3838 (.out1(R3839), .clock(clock), .in1(R3838));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4071 (.out1(R4072), .clock(clock), .in1(R4071));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4249 (.out1(R4250), .clock(clock), .in1(R4249));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4423 (.out1(R4424), .clock(clock), .in1(R4423));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4642 (.out1(R4643), .clock(clock), .in1(R4642));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4806 (.out1(R4807), .clock(clock), .in1(R4806));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4966 (.out1(R4967), .clock(clock), .in1(R4966));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5171 (.out1(R5172), .clock(clock), .in1(R5171));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5321 (.out1(R5322), .clock(clock), .in1(R5321));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5467 (.out1(R5468), .clock(clock), .in1(R5467));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5658 (.out1(R5659), .clock(clock), .in1(R5658));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5794 (.out1(R5795), .clock(clock), .in1(R5794));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5926 (.out1(R5927), .clock(clock), .in1(R5926));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6102 (.out1(R6103), .clock(clock), .in1(R6102));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6223 (.out1(R6224), .clock(clock), .in1(R6223));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6340 (.out1(R6341), .clock(clock), .in1(R6340));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6503 (.out1(R6504), .clock(clock), .in1(R6503));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6610 (.out1(R6611), .clock(clock), .in1(R6610));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6713 (.out1(R6714), .clock(clock), .in1(R6713));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6861 (.out1(R6862), .clock(clock), .in1(R6861));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6954 (.out1(R6955), .clock(clock), .in1(R6954));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7043 (.out1(R7044), .clock(clock), .in1(R7043));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7177 (.out1(R7178), .clock(clock), .in1(R7177));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7256 (.out1(R7257), .clock(clock), .in1(R7256));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7331 (.out1(R7332), .clock(clock), .in1(R7331));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7418 (.out1(R7419), .clock(clock), .in1(_861));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7419 (.out1(R7420), .clock(clock), .in1(_803));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7420 (.out1(R7421), .clock(clock), .in1(_854));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7421 (.out1(R7422), .clock(clock), .in1(_844));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7422 (.out1(R7423), .clock(clock), .in1(_838));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7423 (.out1(R7424), .clock(clock), .in1(_826));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7424 (.out1(R7425), .clock(clock), .in1(_820));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7425 (.out1(R7426), .clock(clock), .in1(_810));
  SRAM op903 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_855),.ADR(R7421));
  SRAM op893 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_845),.ADR(R7422));
  SRAM op887 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_839),.ADR(R7423));
  SRAM op875 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_827),.ADR(R7424));
  SRAM op869 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_821),.ADR(R7425));
  SRAM op859 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_811),.ADR(R7426));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op910 (.out1(_862), .in1(7 'd 64), .in2(R7257));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op852 (.out1(_804), .in1(c88_bitmap_2619_D), .in2(R7420));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op911 (.out1(_863), .in1(R7419), .in2(_862));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op904 (.out1(_856), .in1(7 'd 64), .in2(R7257));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op894 (.out1(_846), .in1(7 'd 64), .in2(R7257));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op876 (.out1(_828), .in1(7 'd 64), .in2(R7257));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2804 (.out1(R2805), .clock(clock), .in1(R2804));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3010 (.out1(R3011), .clock(clock), .in1(R3010));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3212 (.out1(R3213), .clock(clock), .in1(R3212));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3459 (.out1(R3460), .clock(clock), .in1(R3459));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3651 (.out1(R3652), .clock(clock), .in1(R3651));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3839 (.out1(R3840), .clock(clock), .in1(R3839));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4072 (.out1(R4073), .clock(clock), .in1(R4072));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4250 (.out1(R4251), .clock(clock), .in1(R4250));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4424 (.out1(R4425), .clock(clock), .in1(R4424));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4643 (.out1(R4644), .clock(clock), .in1(R4643));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4807 (.out1(R4808), .clock(clock), .in1(R4807));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4967 (.out1(R4968), .clock(clock), .in1(R4967));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5172 (.out1(R5173), .clock(clock), .in1(R5172));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5322 (.out1(R5323), .clock(clock), .in1(R5322));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5468 (.out1(R5469), .clock(clock), .in1(R5468));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5659 (.out1(R5660), .clock(clock), .in1(R5659));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5795 (.out1(R5796), .clock(clock), .in1(R5795));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5927 (.out1(R5928), .clock(clock), .in1(R5927));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6103 (.out1(R6104), .clock(clock), .in1(R6103));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6224 (.out1(R6225), .clock(clock), .in1(R6224));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6341 (.out1(R6342), .clock(clock), .in1(R6341));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6504 (.out1(R6505), .clock(clock), .in1(R6504));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6611 (.out1(R6612), .clock(clock), .in1(R6611));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6714 (.out1(R6715), .clock(clock), .in1(R6714));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6862 (.out1(R6863), .clock(clock), .in1(R6862));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6955 (.out1(R6956), .clock(clock), .in1(R6955));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7044 (.out1(R7045), .clock(clock), .in1(R7044));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7178 (.out1(R7179), .clock(clock), .in1(R7178));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7257 (.out1(R7258), .clock(clock), .in1(R7257));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7332 (.out1(R7333), .clock(clock), .in1(R7332));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7426 (.out1(R7427), .clock(clock), .in1(_855));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7427 (.out1(R7428), .clock(clock), .in1(_845));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7428 (.out1(R7429), .clock(clock), .in1(_839));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7429 (.out1(R7430), .clock(clock), .in1(_827));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7430 (.out1(R7431), .clock(clock), .in1(_821));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7431 (.out1(R7432), .clock(clock), .in1(_811));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7432 (.out1(R7433), .clock(clock), .in1(_804));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7433 (.out1(R7434), .clock(clock), .in1(_863));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7434 (.out1(R7435), .clock(clock), .in1(_856));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7435 (.out1(R7436), .clock(clock), .in1(_846));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7436 (.out1(R7437), .clock(clock), .in1(_828));
  SRAM op853 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_805),.ADR(R7433));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op912 (.out1(_864), .in1(R7434), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op905 (.out1(_857), .in1(R7427), .in2(R7435));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op895 (.out1(_847), .in1(R7428), .in2(R7436));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op888 (.out1(_840), .in1(7 'd 64), .in2(R7258));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op877 (.out1(_829), .in1(R7430), .in2(R7437));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op870 (.out1(_822), .in1(7 'd 64), .in2(R7258));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op860 (.out1(_812), .in1(7 'd 64), .in2(R7258));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op913 (.out1(_865), .in1(_864), .in2(63 'd 6148914691236517205));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op914 (.out1(_866), .in1(_857), .in2(_865));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op896 (.out1(_848), .in1(_847), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op889 (.out1(_841), .in1(R7429), .in2(_840));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op878 (.out1(_830), .in1(_829), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op871 (.out1(_823), .in1(R7431), .in2(_822));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op861 (.out1(_813), .in1(R7432), .in2(_812));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op854 (.out1(_806), .in1(7 'd 64), .in2(R7258));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2805 (.out1(R2806), .clock(clock), .in1(R2805));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3011 (.out1(R3012), .clock(clock), .in1(R3011));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3213 (.out1(R3214), .clock(clock), .in1(R3213));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3460 (.out1(R3461), .clock(clock), .in1(R3460));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3652 (.out1(R3653), .clock(clock), .in1(R3652));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3840 (.out1(R3841), .clock(clock), .in1(R3840));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4073 (.out1(R4074), .clock(clock), .in1(R4073));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4251 (.out1(R4252), .clock(clock), .in1(R4251));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4425 (.out1(R4426), .clock(clock), .in1(R4425));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4644 (.out1(R4645), .clock(clock), .in1(R4644));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4808 (.out1(R4809), .clock(clock), .in1(R4808));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4968 (.out1(R4969), .clock(clock), .in1(R4968));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5173 (.out1(R5174), .clock(clock), .in1(R5173));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5323 (.out1(R5324), .clock(clock), .in1(R5323));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5469 (.out1(R5470), .clock(clock), .in1(R5469));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5660 (.out1(R5661), .clock(clock), .in1(R5660));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5796 (.out1(R5797), .clock(clock), .in1(R5796));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5928 (.out1(R5929), .clock(clock), .in1(R5928));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6104 (.out1(R6105), .clock(clock), .in1(R6104));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6225 (.out1(R6226), .clock(clock), .in1(R6225));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6342 (.out1(R6343), .clock(clock), .in1(R6342));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6505 (.out1(R6506), .clock(clock), .in1(R6505));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6612 (.out1(R6613), .clock(clock), .in1(R6612));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6715 (.out1(R6716), .clock(clock), .in1(R6715));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6863 (.out1(R6864), .clock(clock), .in1(R6863));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6956 (.out1(R6957), .clock(clock), .in1(R6956));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7045 (.out1(R7046), .clock(clock), .in1(R7045));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7179 (.out1(R7180), .clock(clock), .in1(R7179));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7258 (.out1(R7259), .clock(clock), .in1(R7258));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7333 (.out1(R7334), .clock(clock), .in1(R7333));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7437 (.out1(R7438), .clock(clock), .in1(_805));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7438 (.out1(R7439), .clock(clock), .in1(_866));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7439 (.out1(R7440), .clock(clock), .in1(_848));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7440 (.out1(R7441), .clock(clock), .in1(_841));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7441 (.out1(R7442), .clock(clock), .in1(_830));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7442 (.out1(R7443), .clock(clock), .in1(_823));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7443 (.out1(R7444), .clock(clock), .in1(_813));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7444 (.out1(R7445), .clock(clock), .in1(_806));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op846 (.out1(_798), .in1(R7180));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op897 (.out1(_849), .in1(R7440), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op915 (.out1(_867), .in1(R7439), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op898 (.out1(_850), .in1(R7441), .in2(_849));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op879 (.out1(_831), .in1(R7442), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op862 (.out1(_814), .in1(R7444), .in2(1 'd 1));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op880 (.out1(_832), .in1(R7443), .in2(_831));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op855 (.out1(_807), .in1(R7438), .in2(R7445));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op847 (.out1(_799), .in1(_798), .in2(2 'd 2));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op916 (.out1(_868), .in1(_867), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op899 (.out1(_851), .in1(_850), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op863 (.out1(_815), .in1(_814), .in2(63 'd 6148914691236517205));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op917 (.out1(_869), .in1(_851), .in2(_868));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op881 (.out1(_833), .in1(_832), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op864 (.out1(_816), .in1(_807), .in2(_815));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2806 (.out1(R2807), .clock(clock), .in1(R2806));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3012 (.out1(R3013), .clock(clock), .in1(R3012));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3214 (.out1(R3215), .clock(clock), .in1(R3214));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3461 (.out1(R3462), .clock(clock), .in1(R3461));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3653 (.out1(R3654), .clock(clock), .in1(R3653));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3841 (.out1(R3842), .clock(clock), .in1(R3841));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4074 (.out1(R4075), .clock(clock), .in1(R4074));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4252 (.out1(R4253), .clock(clock), .in1(R4252));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4426 (.out1(R4427), .clock(clock), .in1(R4426));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4645 (.out1(R4646), .clock(clock), .in1(R4645));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4809 (.out1(R4810), .clock(clock), .in1(R4809));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4969 (.out1(R4970), .clock(clock), .in1(R4969));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5174 (.out1(R5175), .clock(clock), .in1(R5174));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5324 (.out1(R5325), .clock(clock), .in1(R5324));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5470 (.out1(R5471), .clock(clock), .in1(R5470));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5661 (.out1(R5662), .clock(clock), .in1(R5661));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5797 (.out1(R5798), .clock(clock), .in1(R5797));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5929 (.out1(R5930), .clock(clock), .in1(R5929));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6105 (.out1(R6106), .clock(clock), .in1(R6105));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6226 (.out1(R6227), .clock(clock), .in1(R6226));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6343 (.out1(R6344), .clock(clock), .in1(R6343));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6506 (.out1(R6507), .clock(clock), .in1(R6506));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6613 (.out1(R6614), .clock(clock), .in1(R6613));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6716 (.out1(R6717), .clock(clock), .in1(R6716));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6864 (.out1(R6865), .clock(clock), .in1(R6864));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6957 (.out1(R6958), .clock(clock), .in1(R6957));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7046 (.out1(R7047), .clock(clock), .in1(R7046));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7180 (.out1(R7181), .clock(clock), .in1(R7180));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7259 (.out1(R7260), .clock(clock), .in1(R7259));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7334 (.out1(R7335), .clock(clock), .in1(R7334));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7445 (.out1(R7446), .clock(clock), .in1(_799));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7446 (.out1(R7447), .clock(clock), .in1(_869));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7447 (.out1(R7448), .clock(clock), .in1(_833));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7448 (.out1(R7449), .clock(clock), .in1(_816));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op882 (.out1(_834), .in1(R7448), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op865 (.out1(_817), .in1(R7449), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op918 (.out1(_870), .in1(R7447), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op883 (.out1(_835), .in1(_817), .in2(_834));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op848 (.out1(_800), .in1(c88_popcnt_2624_D), .in2(R7446));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op919 (.out1(_871), .in1(_835), .in2(_870));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op920 (.out1(_872), .in1(_871), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2807 (.out1(R2808), .clock(clock), .in1(R2807));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3013 (.out1(R3014), .clock(clock), .in1(R3013));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3215 (.out1(R3216), .clock(clock), .in1(R3215));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3462 (.out1(R3463), .clock(clock), .in1(R3462));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3654 (.out1(R3655), .clock(clock), .in1(R3654));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3842 (.out1(R3843), .clock(clock), .in1(R3842));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4075 (.out1(R4076), .clock(clock), .in1(R4075));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4253 (.out1(R4254), .clock(clock), .in1(R4253));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4427 (.out1(R4428), .clock(clock), .in1(R4427));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4646 (.out1(R4647), .clock(clock), .in1(R4646));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4810 (.out1(R4811), .clock(clock), .in1(R4810));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4970 (.out1(R4971), .clock(clock), .in1(R4970));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5175 (.out1(R5176), .clock(clock), .in1(R5175));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5325 (.out1(R5326), .clock(clock), .in1(R5325));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5471 (.out1(R5472), .clock(clock), .in1(R5471));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5662 (.out1(R5663), .clock(clock), .in1(R5662));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5798 (.out1(R5799), .clock(clock), .in1(R5798));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5930 (.out1(R5931), .clock(clock), .in1(R5930));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6106 (.out1(R6107), .clock(clock), .in1(R6106));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6227 (.out1(R6228), .clock(clock), .in1(R6227));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6344 (.out1(R6345), .clock(clock), .in1(R6344));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6507 (.out1(R6508), .clock(clock), .in1(R6507));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6614 (.out1(R6615), .clock(clock), .in1(R6614));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6717 (.out1(R6718), .clock(clock), .in1(R6717));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6865 (.out1(R6866), .clock(clock), .in1(R6865));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6958 (.out1(R6959), .clock(clock), .in1(R6958));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7047 (.out1(R7048), .clock(clock), .in1(R7047));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7181 (.out1(R7182), .clock(clock), .in1(R7181));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7260 (.out1(R7261), .clock(clock), .in1(R7260));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7335 (.out1(R7336), .clock(clock), .in1(R7335));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7449 (.out1(R7450), .clock(clock), .in1(_800));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7450 (.out1(R7451), .clock(clock), .in1(_872));
  SRAM op849 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_801),.ADR(R7450));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op921 (.out1(_873), .in1(R7451), .in2(57 'd 72340172838076673));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2808 (.out1(R2809), .clock(clock), .in1(R2808));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3014 (.out1(R3015), .clock(clock), .in1(R3014));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3216 (.out1(R3217), .clock(clock), .in1(R3216));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3463 (.out1(R3464), .clock(clock), .in1(R3463));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3655 (.out1(R3656), .clock(clock), .in1(R3655));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3843 (.out1(R3844), .clock(clock), .in1(R3843));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4076 (.out1(R4077), .clock(clock), .in1(R4076));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4254 (.out1(R4255), .clock(clock), .in1(R4254));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4428 (.out1(R4429), .clock(clock), .in1(R4428));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4647 (.out1(R4648), .clock(clock), .in1(R4647));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4811 (.out1(R4812), .clock(clock), .in1(R4811));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4971 (.out1(R4972), .clock(clock), .in1(R4971));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5176 (.out1(R5177), .clock(clock), .in1(R5176));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5326 (.out1(R5327), .clock(clock), .in1(R5326));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5472 (.out1(R5473), .clock(clock), .in1(R5472));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5663 (.out1(R5664), .clock(clock), .in1(R5663));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5799 (.out1(R5800), .clock(clock), .in1(R5799));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5931 (.out1(R5932), .clock(clock), .in1(R5931));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6107 (.out1(R6108), .clock(clock), .in1(R6107));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6228 (.out1(R6229), .clock(clock), .in1(R6228));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6345 (.out1(R6346), .clock(clock), .in1(R6345));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6508 (.out1(R6509), .clock(clock), .in1(R6508));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6615 (.out1(R6616), .clock(clock), .in1(R6615));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6718 (.out1(R6719), .clock(clock), .in1(R6718));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6866 (.out1(R6867), .clock(clock), .in1(R6866));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6959 (.out1(R6960), .clock(clock), .in1(R6959));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7048 (.out1(R7049), .clock(clock), .in1(R7048));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7182 (.out1(R7183), .clock(clock), .in1(R7182));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7261 (.out1(R7262), .clock(clock), .in1(R7261));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7336 (.out1(R7337), .clock(clock), .in1(R7336));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7451 (.out1(R7452), .clock(clock), .in1(_801));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7452 (.out1(R7453), .clock(clock), .in1(_873));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op922 (.out1(_874), .in1(R7453), .in2(6 'd 56));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op923 (.out1(_875), .in1(_874));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op924 (.out1(ck_idx_2625), .in1(R7452), .in2(_875));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2809 (.out1(R2810), .clock(clock), .in1(R2809));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3015 (.out1(R3016), .clock(clock), .in1(R3015));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3217 (.out1(R3218), .clock(clock), .in1(R3217));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3464 (.out1(R3465), .clock(clock), .in1(R3464));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3656 (.out1(R3657), .clock(clock), .in1(R3656));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3844 (.out1(R3845), .clock(clock), .in1(R3844));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4077 (.out1(R4078), .clock(clock), .in1(R4077));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4255 (.out1(R4256), .clock(clock), .in1(R4255));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4429 (.out1(R4430), .clock(clock), .in1(R4429));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4648 (.out1(R4649), .clock(clock), .in1(R4648));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4812 (.out1(R4813), .clock(clock), .in1(R4812));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4972 (.out1(R4973), .clock(clock), .in1(R4972));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5177 (.out1(R5178), .clock(clock), .in1(R5177));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5327 (.out1(R5328), .clock(clock), .in1(R5327));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5473 (.out1(R5474), .clock(clock), .in1(R5473));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5664 (.out1(R5665), .clock(clock), .in1(R5664));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5800 (.out1(R5801), .clock(clock), .in1(R5800));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5932 (.out1(R5933), .clock(clock), .in1(R5932));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6108 (.out1(R6109), .clock(clock), .in1(R6108));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6229 (.out1(R6230), .clock(clock), .in1(R6229));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6346 (.out1(R6347), .clock(clock), .in1(R6346));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6509 (.out1(R6510), .clock(clock), .in1(R6509));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6616 (.out1(R6617), .clock(clock), .in1(R6616));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6719 (.out1(R6720), .clock(clock), .in1(R6719));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6867 (.out1(R6868), .clock(clock), .in1(R6867));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6960 (.out1(R6961), .clock(clock), .in1(R6960));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7049 (.out1(R7050), .clock(clock), .in1(R7049));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7183 (.out1(R7184), .clock(clock), .in1(R7183));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7262 (.out1(R7263), .clock(clock), .in1(R7262));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7337 (.out1(R7338), .clock(clock), .in1(R7337));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7453 (.out1(R7454), .clock(clock), .in1(ck_idx_2625));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(4), .BITSIZE_out1(32), .PRECISION(32)) op925 (.out1(_876), .in1(R7454), .in2(4 'd 8));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op926 (.out1(_877), .in1(ip2_2595_D), .in2(6 'd 32));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2810 (.out1(R2811), .clock(clock), .in1(R2810));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3016 (.out1(R3017), .clock(clock), .in1(R3016));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3218 (.out1(R3219), .clock(clock), .in1(R3218));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3465 (.out1(R3466), .clock(clock), .in1(R3465));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3657 (.out1(R3658), .clock(clock), .in1(R3657));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3845 (.out1(R3846), .clock(clock), .in1(R3845));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4078 (.out1(R4079), .clock(clock), .in1(R4078));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4256 (.out1(R4257), .clock(clock), .in1(R4256));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4430 (.out1(R4431), .clock(clock), .in1(R4430));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4649 (.out1(R4650), .clock(clock), .in1(R4649));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4813 (.out1(R4814), .clock(clock), .in1(R4813));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4973 (.out1(R4974), .clock(clock), .in1(R4973));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5178 (.out1(R5179), .clock(clock), .in1(R5178));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5328 (.out1(R5329), .clock(clock), .in1(R5328));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5474 (.out1(R5475), .clock(clock), .in1(R5474));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5665 (.out1(R5666), .clock(clock), .in1(R5665));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5801 (.out1(R5802), .clock(clock), .in1(R5801));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5933 (.out1(R5934), .clock(clock), .in1(R5933));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6109 (.out1(R6110), .clock(clock), .in1(R6109));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6230 (.out1(R6231), .clock(clock), .in1(R6230));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6347 (.out1(R6348), .clock(clock), .in1(R6347));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6510 (.out1(R6511), .clock(clock), .in1(R6510));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6617 (.out1(R6618), .clock(clock), .in1(R6617));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6720 (.out1(R6721), .clock(clock), .in1(R6720));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6868 (.out1(R6869), .clock(clock), .in1(R6868));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6961 (.out1(R6962), .clock(clock), .in1(R6961));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7050 (.out1(R7051), .clock(clock), .in1(R7050));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7184 (.out1(R7185), .clock(clock), .in1(R7184));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7263 (.out1(R7264), .clock(clock), .in1(R7263));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7338 (.out1(R7339), .clock(clock), .in1(R7338));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7454 (.out1(R7455), .clock(clock), .in1(_876));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7455 (.out1(R7456), .clock(clock), .in1(_877));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op927 (.out1(_878), .in1(R7456));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(8), .BITSIZE_out1(32)) op928 (.out1(_879), .in1(_878), .in2(8 'd 255));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op929 (.out1(idx_sail_2626), .in1(R7455), .in2(_879));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(3), .BITSIZE_out1(32), .PRECISION(32)) op930 (.out1(idx_2627), .in1(idx_sail_2626), .in2(3 'd 6));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2811 (.out1(R2812), .clock(clock), .in1(R2811));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3017 (.out1(R3018), .clock(clock), .in1(R3017));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3219 (.out1(R3220), .clock(clock), .in1(R3219));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3466 (.out1(R3467), .clock(clock), .in1(R3466));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3658 (.out1(R3659), .clock(clock), .in1(R3658));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3846 (.out1(R3847), .clock(clock), .in1(R3846));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4079 (.out1(R4080), .clock(clock), .in1(R4079));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4257 (.out1(R4258), .clock(clock), .in1(R4257));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4431 (.out1(R4432), .clock(clock), .in1(R4431));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4650 (.out1(R4651), .clock(clock), .in1(R4650));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4814 (.out1(R4815), .clock(clock), .in1(R4814));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4974 (.out1(R4975), .clock(clock), .in1(R4974));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5179 (.out1(R5180), .clock(clock), .in1(R5179));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5329 (.out1(R5330), .clock(clock), .in1(R5329));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5475 (.out1(R5476), .clock(clock), .in1(R5475));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5666 (.out1(R5667), .clock(clock), .in1(R5666));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5802 (.out1(R5803), .clock(clock), .in1(R5802));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5934 (.out1(R5935), .clock(clock), .in1(R5934));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6110 (.out1(R6111), .clock(clock), .in1(R6110));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6231 (.out1(R6232), .clock(clock), .in1(R6231));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6348 (.out1(R6349), .clock(clock), .in1(R6348));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6511 (.out1(R6512), .clock(clock), .in1(R6511));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6618 (.out1(R6619), .clock(clock), .in1(R6618));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6721 (.out1(R6722), .clock(clock), .in1(R6721));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6869 (.out1(R6870), .clock(clock), .in1(R6869));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6962 (.out1(R6963), .clock(clock), .in1(R6962));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7051 (.out1(R7052), .clock(clock), .in1(R7051));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7185 (.out1(R7186), .clock(clock), .in1(R7185));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7264 (.out1(R7265), .clock(clock), .in1(R7264));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7339 (.out1(R7340), .clock(clock), .in1(R7339));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7456 (.out1(R7457), .clock(clock), .in1(idx_sail_2626));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7459 (.out1(R7460), .clock(clock), .in1(idx_2627));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op932 (.out1(_880), .in1(R7460));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op933 (.out1(_881), .in1(_880), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2812 (.out1(R2813), .clock(clock), .in1(R2812));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3018 (.out1(R3019), .clock(clock), .in1(R3018));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3220 (.out1(R3221), .clock(clock), .in1(R3220));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3467 (.out1(R3468), .clock(clock), .in1(R3467));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3659 (.out1(R3660), .clock(clock), .in1(R3659));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3847 (.out1(R3848), .clock(clock), .in1(R3847));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4080 (.out1(R4081), .clock(clock), .in1(R4080));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4258 (.out1(R4259), .clock(clock), .in1(R4258));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4432 (.out1(R4433), .clock(clock), .in1(R4432));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4651 (.out1(R4652), .clock(clock), .in1(R4651));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4815 (.out1(R4816), .clock(clock), .in1(R4815));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4975 (.out1(R4976), .clock(clock), .in1(R4975));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5180 (.out1(R5181), .clock(clock), .in1(R5180));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5330 (.out1(R5331), .clock(clock), .in1(R5330));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5476 (.out1(R5477), .clock(clock), .in1(R5476));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5667 (.out1(R5668), .clock(clock), .in1(R5667));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5803 (.out1(R5804), .clock(clock), .in1(R5803));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5935 (.out1(R5936), .clock(clock), .in1(R5935));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6111 (.out1(R6112), .clock(clock), .in1(R6111));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6232 (.out1(R6233), .clock(clock), .in1(R6232));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6349 (.out1(R6350), .clock(clock), .in1(R6349));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6512 (.out1(R6513), .clock(clock), .in1(R6512));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6619 (.out1(R6620), .clock(clock), .in1(R6619));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6722 (.out1(R6723), .clock(clock), .in1(R6722));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6870 (.out1(R6871), .clock(clock), .in1(R6870));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6963 (.out1(R6964), .clock(clock), .in1(R6963));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7052 (.out1(R7053), .clock(clock), .in1(R7052));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7186 (.out1(R7187), .clock(clock), .in1(R7186));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7265 (.out1(R7266), .clock(clock), .in1(R7265));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7340 (.out1(R7341), .clock(clock), .in1(R7340));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7457 (.out1(R7458), .clock(clock), .in1(R7457));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7460 (.out1(R7461), .clock(clock), .in1(R7460));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7524 (.out1(R7525), .clock(clock), .in1(_881));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op934 (.out1(_882), .in1(c96_bitmap_2629_D), .in2(R7525));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2813 (.out1(R2814), .clock(clock), .in1(R2813));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3019 (.out1(R3020), .clock(clock), .in1(R3019));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3221 (.out1(R3222), .clock(clock), .in1(R3221));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3468 (.out1(R3469), .clock(clock), .in1(R3468));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3660 (.out1(R3661), .clock(clock), .in1(R3660));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3848 (.out1(R3849), .clock(clock), .in1(R3848));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4081 (.out1(R4082), .clock(clock), .in1(R4081));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4259 (.out1(R4260), .clock(clock), .in1(R4259));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4433 (.out1(R4434), .clock(clock), .in1(R4433));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4652 (.out1(R4653), .clock(clock), .in1(R4652));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4816 (.out1(R4817), .clock(clock), .in1(R4816));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4976 (.out1(R4977), .clock(clock), .in1(R4976));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5181 (.out1(R5182), .clock(clock), .in1(R5181));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5331 (.out1(R5332), .clock(clock), .in1(R5331));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5477 (.out1(R5478), .clock(clock), .in1(R5477));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5668 (.out1(R5669), .clock(clock), .in1(R5668));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5804 (.out1(R5805), .clock(clock), .in1(R5804));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5936 (.out1(R5937), .clock(clock), .in1(R5936));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6112 (.out1(R6113), .clock(clock), .in1(R6112));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6233 (.out1(R6234), .clock(clock), .in1(R6233));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6350 (.out1(R6351), .clock(clock), .in1(R6350));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6513 (.out1(R6514), .clock(clock), .in1(R6513));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6620 (.out1(R6621), .clock(clock), .in1(R6620));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6723 (.out1(R6724), .clock(clock), .in1(R6723));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6871 (.out1(R6872), .clock(clock), .in1(R6871));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6964 (.out1(R6965), .clock(clock), .in1(R6964));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7053 (.out1(R7054), .clock(clock), .in1(R7053));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7187 (.out1(R7188), .clock(clock), .in1(R7187));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7266 (.out1(R7267), .clock(clock), .in1(R7266));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7341 (.out1(R7342), .clock(clock), .in1(R7341));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7458 (.out1(R7459), .clock(clock), .in1(R7458));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7461 (.out1(R7462), .clock(clock), .in1(R7461));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7525 (.out1(R7526), .clock(clock), .in1(_882));
  SRAM op935 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_883),.ADR(R7526));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op931 (.out1(off_2628), .in1(R7459), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op936 (.out1(_884), .in1(64 'd 9223372036854775808), .in2(off_2628));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2814 (.out1(R2815), .clock(clock), .in1(R2814));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3020 (.out1(R3021), .clock(clock), .in1(R3020));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3222 (.out1(R3223), .clock(clock), .in1(R3222));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3469 (.out1(R3470), .clock(clock), .in1(R3469));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3661 (.out1(R3662), .clock(clock), .in1(R3661));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3849 (.out1(R3850), .clock(clock), .in1(R3849));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4082 (.out1(R4083), .clock(clock), .in1(R4082));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4260 (.out1(R4261), .clock(clock), .in1(R4260));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4434 (.out1(R4435), .clock(clock), .in1(R4434));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4653 (.out1(R4654), .clock(clock), .in1(R4653));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4817 (.out1(R4818), .clock(clock), .in1(R4817));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4977 (.out1(R4978), .clock(clock), .in1(R4977));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5182 (.out1(R5183), .clock(clock), .in1(R5182));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5332 (.out1(R5333), .clock(clock), .in1(R5332));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5478 (.out1(R5479), .clock(clock), .in1(R5478));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5669 (.out1(R5670), .clock(clock), .in1(R5669));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5805 (.out1(R5806), .clock(clock), .in1(R5805));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5937 (.out1(R5938), .clock(clock), .in1(R5937));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6113 (.out1(R6114), .clock(clock), .in1(R6113));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6234 (.out1(R6235), .clock(clock), .in1(R6234));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6351 (.out1(R6352), .clock(clock), .in1(R6351));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6514 (.out1(R6515), .clock(clock), .in1(R6514));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6621 (.out1(R6622), .clock(clock), .in1(R6621));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6724 (.out1(R6725), .clock(clock), .in1(R6724));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6872 (.out1(R6873), .clock(clock), .in1(R6872));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6965 (.out1(R6966), .clock(clock), .in1(R6965));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7054 (.out1(R7055), .clock(clock), .in1(R7054));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7188 (.out1(R7189), .clock(clock), .in1(R7188));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7267 (.out1(R7268), .clock(clock), .in1(R7267));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7342 (.out1(R7343), .clock(clock), .in1(R7342));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7462 (.out1(R7463), .clock(clock), .in1(R7462));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7526 (.out1(R7527), .clock(clock), .in1(_883));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7527 (.out1(R7528), .clock(clock), .in1(off_2628));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7588 (.out1(R7589), .clock(clock), .in1(_884));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op937 (.out1(_885), .in1(R7527), .in2(R7589));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op938 (.out1(ifout938), .in1(_885), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op999 (.out1(_946), .in1(R7463));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1000 (.out1(_947), .in1(_946), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2815 (.out1(R2816), .clock(clock), .in1(R2815));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3021 (.out1(R3022), .clock(clock), .in1(R3021));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3223 (.out1(R3224), .clock(clock), .in1(R3223));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3470 (.out1(R3471), .clock(clock), .in1(R3470));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3662 (.out1(R3663), .clock(clock), .in1(R3662));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3850 (.out1(R3851), .clock(clock), .in1(R3850));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4083 (.out1(R4084), .clock(clock), .in1(R4083));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4261 (.out1(R4262), .clock(clock), .in1(R4261));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4435 (.out1(R4436), .clock(clock), .in1(R4435));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4654 (.out1(R4655), .clock(clock), .in1(R4654));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4818 (.out1(R4819), .clock(clock), .in1(R4818));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4978 (.out1(R4979), .clock(clock), .in1(R4978));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5183 (.out1(R5184), .clock(clock), .in1(R5183));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5333 (.out1(R5334), .clock(clock), .in1(R5333));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5479 (.out1(R5480), .clock(clock), .in1(R5479));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5670 (.out1(R5671), .clock(clock), .in1(R5670));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5806 (.out1(R5807), .clock(clock), .in1(R5806));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5938 (.out1(R5939), .clock(clock), .in1(R5938));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6114 (.out1(R6115), .clock(clock), .in1(R6114));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6235 (.out1(R6236), .clock(clock), .in1(R6235));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6352 (.out1(R6353), .clock(clock), .in1(R6352));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6515 (.out1(R6516), .clock(clock), .in1(R6515));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6622 (.out1(R6623), .clock(clock), .in1(R6622));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6725 (.out1(R6726), .clock(clock), .in1(R6725));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6873 (.out1(R6874), .clock(clock), .in1(R6873));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6966 (.out1(R6967), .clock(clock), .in1(R6966));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7055 (.out1(R7056), .clock(clock), .in1(R7055));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7189 (.out1(R7190), .clock(clock), .in1(R7189));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7268 (.out1(R7269), .clock(clock), .in1(R7268));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7343 (.out1(R7344), .clock(clock), .in1(R7343));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7463 (.out1(R7464), .clock(clock), .in1(R7463));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7528 (.out1(R7529), .clock(clock), .in1(R7528));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7589 (.out1(R7590), .clock(clock), .in1(ifout938));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7656 (.out1(R7657), .clock(clock), .in1(_947));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op993 (.out1(_940), .in1(R7464));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op983 (.out1(_930), .in1(R7464));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op977 (.out1(_924), .in1(R7464));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op965 (.out1(_912), .in1(R7464));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op959 (.out1(_906), .in1(R7464));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op949 (.out1(_896), .in1(R7464));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op994 (.out1(_941), .in1(_940), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op984 (.out1(_931), .in1(_930), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op978 (.out1(_925), .in1(_924), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op966 (.out1(_913), .in1(_912), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op960 (.out1(_907), .in1(_906), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op950 (.out1(_897), .in1(_896), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1001 (.out1(_948), .in1(c96_bitmap_2629_D), .in2(R7657));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2816 (.out1(R2817), .clock(clock), .in1(R2816));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3022 (.out1(R3023), .clock(clock), .in1(R3022));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3224 (.out1(R3225), .clock(clock), .in1(R3224));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3471 (.out1(R3472), .clock(clock), .in1(R3471));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3663 (.out1(R3664), .clock(clock), .in1(R3663));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3851 (.out1(R3852), .clock(clock), .in1(R3851));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4084 (.out1(R4085), .clock(clock), .in1(R4084));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4262 (.out1(R4263), .clock(clock), .in1(R4262));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4436 (.out1(R4437), .clock(clock), .in1(R4436));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4655 (.out1(R4656), .clock(clock), .in1(R4655));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4819 (.out1(R4820), .clock(clock), .in1(R4819));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4979 (.out1(R4980), .clock(clock), .in1(R4979));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5184 (.out1(R5185), .clock(clock), .in1(R5184));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5334 (.out1(R5335), .clock(clock), .in1(R5334));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5480 (.out1(R5481), .clock(clock), .in1(R5480));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5671 (.out1(R5672), .clock(clock), .in1(R5671));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5807 (.out1(R5808), .clock(clock), .in1(R5807));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5939 (.out1(R5940), .clock(clock), .in1(R5939));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6115 (.out1(R6116), .clock(clock), .in1(R6115));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6236 (.out1(R6237), .clock(clock), .in1(R6236));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6353 (.out1(R6354), .clock(clock), .in1(R6353));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6516 (.out1(R6517), .clock(clock), .in1(R6516));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6623 (.out1(R6624), .clock(clock), .in1(R6623));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6726 (.out1(R6727), .clock(clock), .in1(R6726));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6874 (.out1(R6875), .clock(clock), .in1(R6874));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6967 (.out1(R6968), .clock(clock), .in1(R6967));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7056 (.out1(R7057), .clock(clock), .in1(R7056));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7190 (.out1(R7191), .clock(clock), .in1(R7190));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7269 (.out1(R7270), .clock(clock), .in1(R7269));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7344 (.out1(R7345), .clock(clock), .in1(R7344));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7464 (.out1(R7465), .clock(clock), .in1(R7464));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7529 (.out1(R7530), .clock(clock), .in1(R7529));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7590 (.out1(R7591), .clock(clock), .in1(R7590));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7657 (.out1(R7658), .clock(clock), .in1(_941));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7658 (.out1(R7659), .clock(clock), .in1(_931));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7659 (.out1(R7660), .clock(clock), .in1(_925));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7660 (.out1(R7661), .clock(clock), .in1(_913));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7661 (.out1(R7662), .clock(clock), .in1(_907));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7662 (.out1(R7663), .clock(clock), .in1(_897));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7663 (.out1(R7664), .clock(clock), .in1(_948));
  SRAM op1002 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_949),.ADR(R7664));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op943 (.out1(_890), .in1(R7465));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op944 (.out1(_891), .in1(_890), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op995 (.out1(_942), .in1(c96_bitmap_2629_D), .in2(R7658));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op985 (.out1(_932), .in1(c96_bitmap_2629_D), .in2(R7659));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op979 (.out1(_926), .in1(c96_bitmap_2629_D), .in2(R7660));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op967 (.out1(_914), .in1(c96_bitmap_2629_D), .in2(R7661));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op961 (.out1(_908), .in1(c96_bitmap_2629_D), .in2(R7662));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op951 (.out1(_898), .in1(c96_bitmap_2629_D), .in2(R7663));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2817 (.out1(R2818), .clock(clock), .in1(R2817));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3023 (.out1(R3024), .clock(clock), .in1(R3023));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3225 (.out1(R3226), .clock(clock), .in1(R3225));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3472 (.out1(R3473), .clock(clock), .in1(R3472));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3664 (.out1(R3665), .clock(clock), .in1(R3664));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3852 (.out1(R3853), .clock(clock), .in1(R3852));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4085 (.out1(R4086), .clock(clock), .in1(R4085));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4263 (.out1(R4264), .clock(clock), .in1(R4263));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4437 (.out1(R4438), .clock(clock), .in1(R4437));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4656 (.out1(R4657), .clock(clock), .in1(R4656));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4820 (.out1(R4821), .clock(clock), .in1(R4820));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4980 (.out1(R4981), .clock(clock), .in1(R4980));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5185 (.out1(R5186), .clock(clock), .in1(R5185));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5335 (.out1(R5336), .clock(clock), .in1(R5335));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5481 (.out1(R5482), .clock(clock), .in1(R5481));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5672 (.out1(R5673), .clock(clock), .in1(R5672));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5808 (.out1(R5809), .clock(clock), .in1(R5808));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5940 (.out1(R5941), .clock(clock), .in1(R5940));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6116 (.out1(R6117), .clock(clock), .in1(R6116));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6237 (.out1(R6238), .clock(clock), .in1(R6237));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6354 (.out1(R6355), .clock(clock), .in1(R6354));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6517 (.out1(R6518), .clock(clock), .in1(R6517));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6624 (.out1(R6625), .clock(clock), .in1(R6624));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6727 (.out1(R6728), .clock(clock), .in1(R6727));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6875 (.out1(R6876), .clock(clock), .in1(R6875));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6968 (.out1(R6969), .clock(clock), .in1(R6968));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7057 (.out1(R7058), .clock(clock), .in1(R7057));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7191 (.out1(R7192), .clock(clock), .in1(R7191));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7270 (.out1(R7271), .clock(clock), .in1(R7270));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7345 (.out1(R7346), .clock(clock), .in1(R7345));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7465 (.out1(R7466), .clock(clock), .in1(R7465));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7530 (.out1(R7531), .clock(clock), .in1(R7530));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7591 (.out1(R7592), .clock(clock), .in1(R7591));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7664 (.out1(R7665), .clock(clock), .in1(_949));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7665 (.out1(R7666), .clock(clock), .in1(_891));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7666 (.out1(R7667), .clock(clock), .in1(_942));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7667 (.out1(R7668), .clock(clock), .in1(_932));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7668 (.out1(R7669), .clock(clock), .in1(_926));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7669 (.out1(R7670), .clock(clock), .in1(_914));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7670 (.out1(R7671), .clock(clock), .in1(_908));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7671 (.out1(R7672), .clock(clock), .in1(_898));
  SRAM op996 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_943),.ADR(R7667));
  SRAM op986 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_933),.ADR(R7668));
  SRAM op980 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_927),.ADR(R7669));
  SRAM op968 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_915),.ADR(R7670));
  SRAM op962 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_909),.ADR(R7671));
  SRAM op952 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_899),.ADR(R7672));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1003 (.out1(_950), .in1(7 'd 64), .in2(R7531));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op945 (.out1(_892), .in1(c96_bitmap_2629_D), .in2(R7666));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1004 (.out1(_951), .in1(R7665), .in2(_950));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op997 (.out1(_944), .in1(7 'd 64), .in2(R7531));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op987 (.out1(_934), .in1(7 'd 64), .in2(R7531));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op969 (.out1(_916), .in1(7 'd 64), .in2(R7531));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2818 (.out1(R2819), .clock(clock), .in1(R2818));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3024 (.out1(R3025), .clock(clock), .in1(R3024));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3226 (.out1(R3227), .clock(clock), .in1(R3226));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3473 (.out1(R3474), .clock(clock), .in1(R3473));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3665 (.out1(R3666), .clock(clock), .in1(R3665));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3853 (.out1(R3854), .clock(clock), .in1(R3853));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4086 (.out1(R4087), .clock(clock), .in1(R4086));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4264 (.out1(R4265), .clock(clock), .in1(R4264));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4438 (.out1(R4439), .clock(clock), .in1(R4438));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4657 (.out1(R4658), .clock(clock), .in1(R4657));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4821 (.out1(R4822), .clock(clock), .in1(R4821));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4981 (.out1(R4982), .clock(clock), .in1(R4981));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5186 (.out1(R5187), .clock(clock), .in1(R5186));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5336 (.out1(R5337), .clock(clock), .in1(R5336));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5482 (.out1(R5483), .clock(clock), .in1(R5482));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5673 (.out1(R5674), .clock(clock), .in1(R5673));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5809 (.out1(R5810), .clock(clock), .in1(R5809));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5941 (.out1(R5942), .clock(clock), .in1(R5941));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6117 (.out1(R6118), .clock(clock), .in1(R6117));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6238 (.out1(R6239), .clock(clock), .in1(R6238));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6355 (.out1(R6356), .clock(clock), .in1(R6355));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6518 (.out1(R6519), .clock(clock), .in1(R6518));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6625 (.out1(R6626), .clock(clock), .in1(R6625));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6728 (.out1(R6729), .clock(clock), .in1(R6728));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6876 (.out1(R6877), .clock(clock), .in1(R6876));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6969 (.out1(R6970), .clock(clock), .in1(R6969));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7058 (.out1(R7059), .clock(clock), .in1(R7058));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7192 (.out1(R7193), .clock(clock), .in1(R7192));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7271 (.out1(R7272), .clock(clock), .in1(R7271));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7346 (.out1(R7347), .clock(clock), .in1(R7346));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7466 (.out1(R7467), .clock(clock), .in1(R7466));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7531 (.out1(R7532), .clock(clock), .in1(R7531));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7592 (.out1(R7593), .clock(clock), .in1(R7592));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7672 (.out1(R7673), .clock(clock), .in1(_943));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7673 (.out1(R7674), .clock(clock), .in1(_933));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7674 (.out1(R7675), .clock(clock), .in1(_927));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7675 (.out1(R7676), .clock(clock), .in1(_915));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7676 (.out1(R7677), .clock(clock), .in1(_909));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7677 (.out1(R7678), .clock(clock), .in1(_899));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7678 (.out1(R7679), .clock(clock), .in1(_892));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7679 (.out1(R7680), .clock(clock), .in1(_951));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7680 (.out1(R7681), .clock(clock), .in1(_944));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7681 (.out1(R7682), .clock(clock), .in1(_934));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7682 (.out1(R7683), .clock(clock), .in1(_916));
  SRAM op946 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_893),.ADR(R7679));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1005 (.out1(_952), .in1(R7680), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op998 (.out1(_945), .in1(R7673), .in2(R7681));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op988 (.out1(_935), .in1(R7674), .in2(R7682));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op981 (.out1(_928), .in1(7 'd 64), .in2(R7532));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op970 (.out1(_917), .in1(R7676), .in2(R7683));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op963 (.out1(_910), .in1(7 'd 64), .in2(R7532));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op953 (.out1(_900), .in1(7 'd 64), .in2(R7532));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1006 (.out1(_953), .in1(_952), .in2(63 'd 6148914691236517205));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1007 (.out1(_954), .in1(_945), .in2(_953));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op989 (.out1(_936), .in1(_935), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op982 (.out1(_929), .in1(R7675), .in2(_928));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op971 (.out1(_918), .in1(_917), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op964 (.out1(_911), .in1(R7677), .in2(_910));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op954 (.out1(_901), .in1(R7678), .in2(_900));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op947 (.out1(_894), .in1(7 'd 64), .in2(R7532));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2819 (.out1(R2820), .clock(clock), .in1(R2819));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3025 (.out1(R3026), .clock(clock), .in1(R3025));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3227 (.out1(R3228), .clock(clock), .in1(R3227));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3474 (.out1(R3475), .clock(clock), .in1(R3474));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3666 (.out1(R3667), .clock(clock), .in1(R3666));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3854 (.out1(R3855), .clock(clock), .in1(R3854));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4087 (.out1(R4088), .clock(clock), .in1(R4087));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4265 (.out1(R4266), .clock(clock), .in1(R4265));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4439 (.out1(R4440), .clock(clock), .in1(R4439));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4658 (.out1(R4659), .clock(clock), .in1(R4658));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4822 (.out1(R4823), .clock(clock), .in1(R4822));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4982 (.out1(R4983), .clock(clock), .in1(R4982));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5187 (.out1(R5188), .clock(clock), .in1(R5187));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5337 (.out1(R5338), .clock(clock), .in1(R5337));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5483 (.out1(R5484), .clock(clock), .in1(R5483));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5674 (.out1(R5675), .clock(clock), .in1(R5674));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5810 (.out1(R5811), .clock(clock), .in1(R5810));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5942 (.out1(R5943), .clock(clock), .in1(R5942));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6118 (.out1(R6119), .clock(clock), .in1(R6118));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6239 (.out1(R6240), .clock(clock), .in1(R6239));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6356 (.out1(R6357), .clock(clock), .in1(R6356));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6519 (.out1(R6520), .clock(clock), .in1(R6519));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6626 (.out1(R6627), .clock(clock), .in1(R6626));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6729 (.out1(R6730), .clock(clock), .in1(R6729));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6877 (.out1(R6878), .clock(clock), .in1(R6877));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6970 (.out1(R6971), .clock(clock), .in1(R6970));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7059 (.out1(R7060), .clock(clock), .in1(R7059));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7193 (.out1(R7194), .clock(clock), .in1(R7193));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7272 (.out1(R7273), .clock(clock), .in1(R7272));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7347 (.out1(R7348), .clock(clock), .in1(R7347));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7467 (.out1(R7468), .clock(clock), .in1(R7467));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7532 (.out1(R7533), .clock(clock), .in1(R7532));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7593 (.out1(R7594), .clock(clock), .in1(R7593));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7683 (.out1(R7684), .clock(clock), .in1(_893));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7684 (.out1(R7685), .clock(clock), .in1(_954));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7685 (.out1(R7686), .clock(clock), .in1(_936));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7686 (.out1(R7687), .clock(clock), .in1(_929));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7687 (.out1(R7688), .clock(clock), .in1(_918));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7688 (.out1(R7689), .clock(clock), .in1(_911));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7689 (.out1(R7690), .clock(clock), .in1(_901));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7690 (.out1(R7691), .clock(clock), .in1(_894));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op939 (.out1(_886), .in1(R7468));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op990 (.out1(_937), .in1(R7686), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1008 (.out1(_955), .in1(R7685), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op991 (.out1(_938), .in1(R7687), .in2(_937));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op972 (.out1(_919), .in1(R7688), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op955 (.out1(_902), .in1(R7690), .in2(1 'd 1));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op973 (.out1(_920), .in1(R7689), .in2(_919));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op948 (.out1(_895), .in1(R7684), .in2(R7691));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op940 (.out1(_887), .in1(_886), .in2(2 'd 2));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1009 (.out1(_956), .in1(_955), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op992 (.out1(_939), .in1(_938), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op956 (.out1(_903), .in1(_902), .in2(63 'd 6148914691236517205));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1010 (.out1(_957), .in1(_939), .in2(_956));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op974 (.out1(_921), .in1(_920), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op957 (.out1(_904), .in1(_895), .in2(_903));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2820 (.out1(R2821), .clock(clock), .in1(R2820));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3026 (.out1(R3027), .clock(clock), .in1(R3026));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3228 (.out1(R3229), .clock(clock), .in1(R3228));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3475 (.out1(R3476), .clock(clock), .in1(R3475));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3667 (.out1(R3668), .clock(clock), .in1(R3667));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3855 (.out1(R3856), .clock(clock), .in1(R3855));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4088 (.out1(R4089), .clock(clock), .in1(R4088));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4266 (.out1(R4267), .clock(clock), .in1(R4266));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4440 (.out1(R4441), .clock(clock), .in1(R4440));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4659 (.out1(R4660), .clock(clock), .in1(R4659));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4823 (.out1(R4824), .clock(clock), .in1(R4823));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4983 (.out1(R4984), .clock(clock), .in1(R4983));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5188 (.out1(R5189), .clock(clock), .in1(R5188));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5338 (.out1(R5339), .clock(clock), .in1(R5338));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5484 (.out1(R5485), .clock(clock), .in1(R5484));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5675 (.out1(R5676), .clock(clock), .in1(R5675));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5811 (.out1(R5812), .clock(clock), .in1(R5811));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5943 (.out1(R5944), .clock(clock), .in1(R5943));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6119 (.out1(R6120), .clock(clock), .in1(R6119));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6240 (.out1(R6241), .clock(clock), .in1(R6240));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6357 (.out1(R6358), .clock(clock), .in1(R6357));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6520 (.out1(R6521), .clock(clock), .in1(R6520));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6627 (.out1(R6628), .clock(clock), .in1(R6627));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6730 (.out1(R6731), .clock(clock), .in1(R6730));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6878 (.out1(R6879), .clock(clock), .in1(R6878));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6971 (.out1(R6972), .clock(clock), .in1(R6971));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7060 (.out1(R7061), .clock(clock), .in1(R7060));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7194 (.out1(R7195), .clock(clock), .in1(R7194));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7273 (.out1(R7274), .clock(clock), .in1(R7273));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7348 (.out1(R7349), .clock(clock), .in1(R7348));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7468 (.out1(R7469), .clock(clock), .in1(R7468));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7533 (.out1(R7534), .clock(clock), .in1(R7533));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7594 (.out1(R7595), .clock(clock), .in1(R7594));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7691 (.out1(R7692), .clock(clock), .in1(_887));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7692 (.out1(R7693), .clock(clock), .in1(_957));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7693 (.out1(R7694), .clock(clock), .in1(_921));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7694 (.out1(R7695), .clock(clock), .in1(_904));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op975 (.out1(_922), .in1(R7694), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op958 (.out1(_905), .in1(R7695), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op1011 (.out1(_958), .in1(R7693), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op976 (.out1(_923), .in1(_905), .in2(_922));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op941 (.out1(_888), .in1(c96_popcnt_2634_D), .in2(R7692));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1012 (.out1(_959), .in1(_923), .in2(_958));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op1013 (.out1(_960), .in1(_959), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2821 (.out1(R2822), .clock(clock), .in1(R2821));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3027 (.out1(R3028), .clock(clock), .in1(R3027));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3229 (.out1(R3230), .clock(clock), .in1(R3229));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3476 (.out1(R3477), .clock(clock), .in1(R3476));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3668 (.out1(R3669), .clock(clock), .in1(R3668));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3856 (.out1(R3857), .clock(clock), .in1(R3856));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4089 (.out1(R4090), .clock(clock), .in1(R4089));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4267 (.out1(R4268), .clock(clock), .in1(R4267));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4441 (.out1(R4442), .clock(clock), .in1(R4441));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4660 (.out1(R4661), .clock(clock), .in1(R4660));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4824 (.out1(R4825), .clock(clock), .in1(R4824));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4984 (.out1(R4985), .clock(clock), .in1(R4984));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5189 (.out1(R5190), .clock(clock), .in1(R5189));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5339 (.out1(R5340), .clock(clock), .in1(R5339));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5485 (.out1(R5486), .clock(clock), .in1(R5485));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5676 (.out1(R5677), .clock(clock), .in1(R5676));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5812 (.out1(R5813), .clock(clock), .in1(R5812));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5944 (.out1(R5945), .clock(clock), .in1(R5944));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6120 (.out1(R6121), .clock(clock), .in1(R6120));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6241 (.out1(R6242), .clock(clock), .in1(R6241));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6358 (.out1(R6359), .clock(clock), .in1(R6358));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6521 (.out1(R6522), .clock(clock), .in1(R6521));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6628 (.out1(R6629), .clock(clock), .in1(R6628));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6731 (.out1(R6732), .clock(clock), .in1(R6731));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6879 (.out1(R6880), .clock(clock), .in1(R6879));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6972 (.out1(R6973), .clock(clock), .in1(R6972));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7061 (.out1(R7062), .clock(clock), .in1(R7061));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7195 (.out1(R7196), .clock(clock), .in1(R7195));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7274 (.out1(R7275), .clock(clock), .in1(R7274));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7349 (.out1(R7350), .clock(clock), .in1(R7349));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7469 (.out1(R7470), .clock(clock), .in1(R7469));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7534 (.out1(R7535), .clock(clock), .in1(R7534));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7595 (.out1(R7596), .clock(clock), .in1(R7595));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7695 (.out1(R7696), .clock(clock), .in1(_888));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7696 (.out1(R7697), .clock(clock), .in1(_960));
  SRAM op942 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_889),.ADR(R7696));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op1014 (.out1(_961), .in1(R7697), .in2(57 'd 72340172838076673));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2822 (.out1(R2823), .clock(clock), .in1(R2822));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3028 (.out1(R3029), .clock(clock), .in1(R3028));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3230 (.out1(R3231), .clock(clock), .in1(R3230));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3477 (.out1(R3478), .clock(clock), .in1(R3477));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3669 (.out1(R3670), .clock(clock), .in1(R3669));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3857 (.out1(R3858), .clock(clock), .in1(R3857));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4090 (.out1(R4091), .clock(clock), .in1(R4090));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4268 (.out1(R4269), .clock(clock), .in1(R4268));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4442 (.out1(R4443), .clock(clock), .in1(R4442));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4661 (.out1(R4662), .clock(clock), .in1(R4661));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4825 (.out1(R4826), .clock(clock), .in1(R4825));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4985 (.out1(R4986), .clock(clock), .in1(R4985));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5190 (.out1(R5191), .clock(clock), .in1(R5190));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5340 (.out1(R5341), .clock(clock), .in1(R5340));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5486 (.out1(R5487), .clock(clock), .in1(R5486));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5677 (.out1(R5678), .clock(clock), .in1(R5677));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5813 (.out1(R5814), .clock(clock), .in1(R5813));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5945 (.out1(R5946), .clock(clock), .in1(R5945));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6121 (.out1(R6122), .clock(clock), .in1(R6121));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6242 (.out1(R6243), .clock(clock), .in1(R6242));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6359 (.out1(R6360), .clock(clock), .in1(R6359));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6522 (.out1(R6523), .clock(clock), .in1(R6522));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6629 (.out1(R6630), .clock(clock), .in1(R6629));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6732 (.out1(R6733), .clock(clock), .in1(R6732));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6880 (.out1(R6881), .clock(clock), .in1(R6880));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6973 (.out1(R6974), .clock(clock), .in1(R6973));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7062 (.out1(R7063), .clock(clock), .in1(R7062));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7196 (.out1(R7197), .clock(clock), .in1(R7196));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7275 (.out1(R7276), .clock(clock), .in1(R7275));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7350 (.out1(R7351), .clock(clock), .in1(R7350));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7470 (.out1(R7471), .clock(clock), .in1(R7470));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7535 (.out1(R7536), .clock(clock), .in1(R7535));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7596 (.out1(R7597), .clock(clock), .in1(R7596));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7697 (.out1(R7698), .clock(clock), .in1(_889));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7698 (.out1(R7699), .clock(clock), .in1(_961));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op1015 (.out1(_962), .in1(R7699), .in2(6 'd 56));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1016 (.out1(_963), .in1(_962));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1017 (.out1(ck_idx_2635), .in1(R7698), .in2(_963));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2823 (.out1(R2824), .clock(clock), .in1(R2823));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3029 (.out1(R3030), .clock(clock), .in1(R3029));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3231 (.out1(R3232), .clock(clock), .in1(R3231));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3478 (.out1(R3479), .clock(clock), .in1(R3478));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3670 (.out1(R3671), .clock(clock), .in1(R3670));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3858 (.out1(R3859), .clock(clock), .in1(R3858));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4091 (.out1(R4092), .clock(clock), .in1(R4091));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4269 (.out1(R4270), .clock(clock), .in1(R4269));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4443 (.out1(R4444), .clock(clock), .in1(R4443));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4662 (.out1(R4663), .clock(clock), .in1(R4662));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4826 (.out1(R4827), .clock(clock), .in1(R4826));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4986 (.out1(R4987), .clock(clock), .in1(R4986));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5191 (.out1(R5192), .clock(clock), .in1(R5191));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5341 (.out1(R5342), .clock(clock), .in1(R5341));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5487 (.out1(R5488), .clock(clock), .in1(R5487));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5678 (.out1(R5679), .clock(clock), .in1(R5678));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5814 (.out1(R5815), .clock(clock), .in1(R5814));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5946 (.out1(R5947), .clock(clock), .in1(R5946));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6122 (.out1(R6123), .clock(clock), .in1(R6122));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6243 (.out1(R6244), .clock(clock), .in1(R6243));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6360 (.out1(R6361), .clock(clock), .in1(R6360));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6523 (.out1(R6524), .clock(clock), .in1(R6523));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6630 (.out1(R6631), .clock(clock), .in1(R6630));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6733 (.out1(R6734), .clock(clock), .in1(R6733));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6881 (.out1(R6882), .clock(clock), .in1(R6881));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6974 (.out1(R6975), .clock(clock), .in1(R6974));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7063 (.out1(R7064), .clock(clock), .in1(R7063));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7197 (.out1(R7198), .clock(clock), .in1(R7197));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7276 (.out1(R7277), .clock(clock), .in1(R7276));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7351 (.out1(R7352), .clock(clock), .in1(R7351));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7471 (.out1(R7472), .clock(clock), .in1(R7471));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7536 (.out1(R7537), .clock(clock), .in1(R7536));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7597 (.out1(R7598), .clock(clock), .in1(R7597));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7699 (.out1(R7700), .clock(clock), .in1(ck_idx_2635));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(4), .BITSIZE_out1(32), .PRECISION(32)) op1018 (.out1(_964), .in1(R7700), .in2(4 'd 8));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(5), .BITSIZE_out1(64), .PRECISION(64)) op1019 (.out1(_965), .in1(ip2_2595_D), .in2(5 'd 24));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2824 (.out1(R2825), .clock(clock), .in1(R2824));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3030 (.out1(R3031), .clock(clock), .in1(R3030));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3232 (.out1(R3233), .clock(clock), .in1(R3232));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3479 (.out1(R3480), .clock(clock), .in1(R3479));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3671 (.out1(R3672), .clock(clock), .in1(R3671));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3859 (.out1(R3860), .clock(clock), .in1(R3859));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4092 (.out1(R4093), .clock(clock), .in1(R4092));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4270 (.out1(R4271), .clock(clock), .in1(R4270));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4444 (.out1(R4445), .clock(clock), .in1(R4444));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4663 (.out1(R4664), .clock(clock), .in1(R4663));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4827 (.out1(R4828), .clock(clock), .in1(R4827));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4987 (.out1(R4988), .clock(clock), .in1(R4987));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5192 (.out1(R5193), .clock(clock), .in1(R5192));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5342 (.out1(R5343), .clock(clock), .in1(R5342));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5488 (.out1(R5489), .clock(clock), .in1(R5488));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5679 (.out1(R5680), .clock(clock), .in1(R5679));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5815 (.out1(R5816), .clock(clock), .in1(R5815));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5947 (.out1(R5948), .clock(clock), .in1(R5947));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6123 (.out1(R6124), .clock(clock), .in1(R6123));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6244 (.out1(R6245), .clock(clock), .in1(R6244));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6361 (.out1(R6362), .clock(clock), .in1(R6361));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6524 (.out1(R6525), .clock(clock), .in1(R6524));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6631 (.out1(R6632), .clock(clock), .in1(R6631));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6734 (.out1(R6735), .clock(clock), .in1(R6734));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6882 (.out1(R6883), .clock(clock), .in1(R6882));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6975 (.out1(R6976), .clock(clock), .in1(R6975));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7064 (.out1(R7065), .clock(clock), .in1(R7064));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7198 (.out1(R7199), .clock(clock), .in1(R7198));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7277 (.out1(R7278), .clock(clock), .in1(R7277));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7352 (.out1(R7353), .clock(clock), .in1(R7352));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7472 (.out1(R7473), .clock(clock), .in1(R7472));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7537 (.out1(R7538), .clock(clock), .in1(R7537));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7598 (.out1(R7599), .clock(clock), .in1(R7598));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7700 (.out1(R7701), .clock(clock), .in1(_964));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7701 (.out1(R7702), .clock(clock), .in1(_965));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1020 (.out1(_966), .in1(R7702));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(8), .BITSIZE_out1(32)) op1021 (.out1(_967), .in1(_966), .in2(8 'd 255));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1022 (.out1(idx_sail_2636), .in1(R7701), .in2(_967));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(3), .BITSIZE_out1(32), .PRECISION(32)) op1023 (.out1(idx_2637), .in1(idx_sail_2636), .in2(3 'd 6));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2825 (.out1(R2826), .clock(clock), .in1(R2825));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3031 (.out1(R3032), .clock(clock), .in1(R3031));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3233 (.out1(R3234), .clock(clock), .in1(R3233));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3480 (.out1(R3481), .clock(clock), .in1(R3480));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3672 (.out1(R3673), .clock(clock), .in1(R3672));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3860 (.out1(R3861), .clock(clock), .in1(R3860));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4093 (.out1(R4094), .clock(clock), .in1(R4093));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4271 (.out1(R4272), .clock(clock), .in1(R4271));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4445 (.out1(R4446), .clock(clock), .in1(R4445));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4664 (.out1(R4665), .clock(clock), .in1(R4664));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4828 (.out1(R4829), .clock(clock), .in1(R4828));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4988 (.out1(R4989), .clock(clock), .in1(R4988));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5193 (.out1(R5194), .clock(clock), .in1(R5193));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5343 (.out1(R5344), .clock(clock), .in1(R5343));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5489 (.out1(R5490), .clock(clock), .in1(R5489));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5680 (.out1(R5681), .clock(clock), .in1(R5680));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5816 (.out1(R5817), .clock(clock), .in1(R5816));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5948 (.out1(R5949), .clock(clock), .in1(R5948));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6124 (.out1(R6125), .clock(clock), .in1(R6124));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6245 (.out1(R6246), .clock(clock), .in1(R6245));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6362 (.out1(R6363), .clock(clock), .in1(R6362));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6525 (.out1(R6526), .clock(clock), .in1(R6525));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6632 (.out1(R6633), .clock(clock), .in1(R6632));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6735 (.out1(R6736), .clock(clock), .in1(R6735));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6883 (.out1(R6884), .clock(clock), .in1(R6883));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6976 (.out1(R6977), .clock(clock), .in1(R6976));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7065 (.out1(R7066), .clock(clock), .in1(R7065));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7199 (.out1(R7200), .clock(clock), .in1(R7199));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7278 (.out1(R7279), .clock(clock), .in1(R7278));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7353 (.out1(R7354), .clock(clock), .in1(R7353));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7473 (.out1(R7474), .clock(clock), .in1(R7473));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7538 (.out1(R7539), .clock(clock), .in1(R7538));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7599 (.out1(R7600), .clock(clock), .in1(R7599));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7702 (.out1(R7703), .clock(clock), .in1(idx_sail_2636));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7705 (.out1(R7706), .clock(clock), .in1(idx_2637));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1025 (.out1(_968), .in1(R7706));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1026 (.out1(_969), .in1(_968), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2826 (.out1(R2827), .clock(clock), .in1(R2826));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3032 (.out1(R3033), .clock(clock), .in1(R3032));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3234 (.out1(R3235), .clock(clock), .in1(R3234));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3481 (.out1(R3482), .clock(clock), .in1(R3481));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3673 (.out1(R3674), .clock(clock), .in1(R3673));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3861 (.out1(R3862), .clock(clock), .in1(R3861));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4094 (.out1(R4095), .clock(clock), .in1(R4094));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4272 (.out1(R4273), .clock(clock), .in1(R4272));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4446 (.out1(R4447), .clock(clock), .in1(R4446));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4665 (.out1(R4666), .clock(clock), .in1(R4665));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4829 (.out1(R4830), .clock(clock), .in1(R4829));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4989 (.out1(R4990), .clock(clock), .in1(R4989));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5194 (.out1(R5195), .clock(clock), .in1(R5194));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5344 (.out1(R5345), .clock(clock), .in1(R5344));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5490 (.out1(R5491), .clock(clock), .in1(R5490));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5681 (.out1(R5682), .clock(clock), .in1(R5681));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5817 (.out1(R5818), .clock(clock), .in1(R5817));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5949 (.out1(R5950), .clock(clock), .in1(R5949));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6125 (.out1(R6126), .clock(clock), .in1(R6125));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6246 (.out1(R6247), .clock(clock), .in1(R6246));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6363 (.out1(R6364), .clock(clock), .in1(R6363));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6526 (.out1(R6527), .clock(clock), .in1(R6526));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6633 (.out1(R6634), .clock(clock), .in1(R6633));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6736 (.out1(R6737), .clock(clock), .in1(R6736));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6884 (.out1(R6885), .clock(clock), .in1(R6884));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6977 (.out1(R6978), .clock(clock), .in1(R6977));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7066 (.out1(R7067), .clock(clock), .in1(R7066));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7200 (.out1(R7201), .clock(clock), .in1(R7200));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7279 (.out1(R7280), .clock(clock), .in1(R7279));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7354 (.out1(R7355), .clock(clock), .in1(R7354));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7474 (.out1(R7475), .clock(clock), .in1(R7474));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7539 (.out1(R7540), .clock(clock), .in1(R7539));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7600 (.out1(R7601), .clock(clock), .in1(R7600));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7703 (.out1(R7704), .clock(clock), .in1(R7703));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7706 (.out1(R7707), .clock(clock), .in1(R7706));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7756 (.out1(R7757), .clock(clock), .in1(_969));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1027 (.out1(_970), .in1(c104_bitmap_2639_D), .in2(R7757));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2827 (.out1(R2828), .clock(clock), .in1(R2827));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3033 (.out1(R3034), .clock(clock), .in1(R3033));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3235 (.out1(R3236), .clock(clock), .in1(R3235));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3482 (.out1(R3483), .clock(clock), .in1(R3482));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3674 (.out1(R3675), .clock(clock), .in1(R3674));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3862 (.out1(R3863), .clock(clock), .in1(R3862));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4095 (.out1(R4096), .clock(clock), .in1(R4095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4273 (.out1(R4274), .clock(clock), .in1(R4273));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4447 (.out1(R4448), .clock(clock), .in1(R4447));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4666 (.out1(R4667), .clock(clock), .in1(R4666));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4830 (.out1(R4831), .clock(clock), .in1(R4830));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4990 (.out1(R4991), .clock(clock), .in1(R4990));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5195 (.out1(R5196), .clock(clock), .in1(R5195));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5345 (.out1(R5346), .clock(clock), .in1(R5345));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5491 (.out1(R5492), .clock(clock), .in1(R5491));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5682 (.out1(R5683), .clock(clock), .in1(R5682));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5818 (.out1(R5819), .clock(clock), .in1(R5818));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5950 (.out1(R5951), .clock(clock), .in1(R5950));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6126 (.out1(R6127), .clock(clock), .in1(R6126));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6247 (.out1(R6248), .clock(clock), .in1(R6247));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6364 (.out1(R6365), .clock(clock), .in1(R6364));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6527 (.out1(R6528), .clock(clock), .in1(R6527));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6634 (.out1(R6635), .clock(clock), .in1(R6634));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6737 (.out1(R6738), .clock(clock), .in1(R6737));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6885 (.out1(R6886), .clock(clock), .in1(R6885));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6978 (.out1(R6979), .clock(clock), .in1(R6978));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7067 (.out1(R7068), .clock(clock), .in1(R7067));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7201 (.out1(R7202), .clock(clock), .in1(R7201));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7280 (.out1(R7281), .clock(clock), .in1(R7280));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7355 (.out1(R7356), .clock(clock), .in1(R7355));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7475 (.out1(R7476), .clock(clock), .in1(R7475));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7540 (.out1(R7541), .clock(clock), .in1(R7540));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7601 (.out1(R7602), .clock(clock), .in1(R7601));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7704 (.out1(R7705), .clock(clock), .in1(R7704));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7707 (.out1(R7708), .clock(clock), .in1(R7707));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7757 (.out1(R7758), .clock(clock), .in1(_970));
  SRAM op1028 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_971),.ADR(R7758));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op1024 (.out1(off_2638), .in1(R7705), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1029 (.out1(_972), .in1(64 'd 9223372036854775808), .in2(off_2638));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2828 (.out1(R2829), .clock(clock), .in1(R2828));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3034 (.out1(R3035), .clock(clock), .in1(R3034));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3236 (.out1(R3237), .clock(clock), .in1(R3236));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3483 (.out1(R3484), .clock(clock), .in1(R3483));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3675 (.out1(R3676), .clock(clock), .in1(R3675));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3863 (.out1(R3864), .clock(clock), .in1(R3863));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4096 (.out1(R4097), .clock(clock), .in1(R4096));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4274 (.out1(R4275), .clock(clock), .in1(R4274));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4448 (.out1(R4449), .clock(clock), .in1(R4448));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4667 (.out1(R4668), .clock(clock), .in1(R4667));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4831 (.out1(R4832), .clock(clock), .in1(R4831));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4991 (.out1(R4992), .clock(clock), .in1(R4991));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5196 (.out1(R5197), .clock(clock), .in1(R5196));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5346 (.out1(R5347), .clock(clock), .in1(R5346));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5492 (.out1(R5493), .clock(clock), .in1(R5492));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5683 (.out1(R5684), .clock(clock), .in1(R5683));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5819 (.out1(R5820), .clock(clock), .in1(R5819));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5951 (.out1(R5952), .clock(clock), .in1(R5951));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6127 (.out1(R6128), .clock(clock), .in1(R6127));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6248 (.out1(R6249), .clock(clock), .in1(R6248));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6365 (.out1(R6366), .clock(clock), .in1(R6365));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6528 (.out1(R6529), .clock(clock), .in1(R6528));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6635 (.out1(R6636), .clock(clock), .in1(R6635));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6738 (.out1(R6739), .clock(clock), .in1(R6738));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6886 (.out1(R6887), .clock(clock), .in1(R6886));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6979 (.out1(R6980), .clock(clock), .in1(R6979));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7068 (.out1(R7069), .clock(clock), .in1(R7068));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7202 (.out1(R7203), .clock(clock), .in1(R7202));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7281 (.out1(R7282), .clock(clock), .in1(R7281));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7356 (.out1(R7357), .clock(clock), .in1(R7356));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7476 (.out1(R7477), .clock(clock), .in1(R7476));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7541 (.out1(R7542), .clock(clock), .in1(R7541));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7602 (.out1(R7603), .clock(clock), .in1(R7602));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7708 (.out1(R7709), .clock(clock), .in1(R7708));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7758 (.out1(R7759), .clock(clock), .in1(_971));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7759 (.out1(R7760), .clock(clock), .in1(off_2638));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7806 (.out1(R7807), .clock(clock), .in1(_972));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1030 (.out1(_973), .in1(R7759), .in2(R7807));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op1031 (.out1(ifout1031), .in1(_973), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1092 (.out1(_1034), .in1(R7709));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1093 (.out1(_1035), .in1(_1034), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2829 (.out1(R2830), .clock(clock), .in1(R2829));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3035 (.out1(R3036), .clock(clock), .in1(R3035));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3237 (.out1(R3238), .clock(clock), .in1(R3237));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3484 (.out1(R3485), .clock(clock), .in1(R3484));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3676 (.out1(R3677), .clock(clock), .in1(R3676));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3864 (.out1(R3865), .clock(clock), .in1(R3864));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4097 (.out1(R4098), .clock(clock), .in1(R4097));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4275 (.out1(R4276), .clock(clock), .in1(R4275));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4449 (.out1(R4450), .clock(clock), .in1(R4449));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4668 (.out1(R4669), .clock(clock), .in1(R4668));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4832 (.out1(R4833), .clock(clock), .in1(R4832));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4992 (.out1(R4993), .clock(clock), .in1(R4992));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5197 (.out1(R5198), .clock(clock), .in1(R5197));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5347 (.out1(R5348), .clock(clock), .in1(R5347));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5493 (.out1(R5494), .clock(clock), .in1(R5493));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5684 (.out1(R5685), .clock(clock), .in1(R5684));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5820 (.out1(R5821), .clock(clock), .in1(R5820));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5952 (.out1(R5953), .clock(clock), .in1(R5952));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6128 (.out1(R6129), .clock(clock), .in1(R6128));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6249 (.out1(R6250), .clock(clock), .in1(R6249));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6366 (.out1(R6367), .clock(clock), .in1(R6366));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6529 (.out1(R6530), .clock(clock), .in1(R6529));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6636 (.out1(R6637), .clock(clock), .in1(R6636));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6739 (.out1(R6740), .clock(clock), .in1(R6739));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6887 (.out1(R6888), .clock(clock), .in1(R6887));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6980 (.out1(R6981), .clock(clock), .in1(R6980));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7069 (.out1(R7070), .clock(clock), .in1(R7069));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7203 (.out1(R7204), .clock(clock), .in1(R7203));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7282 (.out1(R7283), .clock(clock), .in1(R7282));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7357 (.out1(R7358), .clock(clock), .in1(R7357));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7477 (.out1(R7478), .clock(clock), .in1(R7477));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7542 (.out1(R7543), .clock(clock), .in1(R7542));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7603 (.out1(R7604), .clock(clock), .in1(R7603));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7709 (.out1(R7710), .clock(clock), .in1(R7709));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7760 (.out1(R7761), .clock(clock), .in1(R7760));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7807 (.out1(R7808), .clock(clock), .in1(ifout1031));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7860 (.out1(R7861), .clock(clock), .in1(_1035));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1086 (.out1(_1028), .in1(R7710));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1076 (.out1(_1018), .in1(R7710));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1070 (.out1(_1012), .in1(R7710));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1058 (.out1(_1000), .in1(R7710));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1052 (.out1(_994), .in1(R7710));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1042 (.out1(_984), .in1(R7710));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1087 (.out1(_1029), .in1(_1028), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1077 (.out1(_1019), .in1(_1018), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1071 (.out1(_1013), .in1(_1012), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1059 (.out1(_1001), .in1(_1000), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1053 (.out1(_995), .in1(_994), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1043 (.out1(_985), .in1(_984), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1094 (.out1(_1036), .in1(c104_bitmap_2639_D), .in2(R7861));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2830 (.out1(R2831), .clock(clock), .in1(R2830));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3036 (.out1(R3037), .clock(clock), .in1(R3036));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3238 (.out1(R3239), .clock(clock), .in1(R3238));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3485 (.out1(R3486), .clock(clock), .in1(R3485));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3677 (.out1(R3678), .clock(clock), .in1(R3677));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3865 (.out1(R3866), .clock(clock), .in1(R3865));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4098 (.out1(R4099), .clock(clock), .in1(R4098));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4276 (.out1(R4277), .clock(clock), .in1(R4276));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4450 (.out1(R4451), .clock(clock), .in1(R4450));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4669 (.out1(R4670), .clock(clock), .in1(R4669));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4833 (.out1(R4834), .clock(clock), .in1(R4833));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4993 (.out1(R4994), .clock(clock), .in1(R4993));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5198 (.out1(R5199), .clock(clock), .in1(R5198));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5348 (.out1(R5349), .clock(clock), .in1(R5348));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5494 (.out1(R5495), .clock(clock), .in1(R5494));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5685 (.out1(R5686), .clock(clock), .in1(R5685));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5821 (.out1(R5822), .clock(clock), .in1(R5821));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5953 (.out1(R5954), .clock(clock), .in1(R5953));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6129 (.out1(R6130), .clock(clock), .in1(R6129));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6250 (.out1(R6251), .clock(clock), .in1(R6250));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6367 (.out1(R6368), .clock(clock), .in1(R6367));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6530 (.out1(R6531), .clock(clock), .in1(R6530));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6637 (.out1(R6638), .clock(clock), .in1(R6637));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6740 (.out1(R6741), .clock(clock), .in1(R6740));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6888 (.out1(R6889), .clock(clock), .in1(R6888));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6981 (.out1(R6982), .clock(clock), .in1(R6981));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7070 (.out1(R7071), .clock(clock), .in1(R7070));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7204 (.out1(R7205), .clock(clock), .in1(R7204));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7283 (.out1(R7284), .clock(clock), .in1(R7283));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7358 (.out1(R7359), .clock(clock), .in1(R7358));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7478 (.out1(R7479), .clock(clock), .in1(R7478));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7543 (.out1(R7544), .clock(clock), .in1(R7543));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7604 (.out1(R7605), .clock(clock), .in1(R7604));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7710 (.out1(R7711), .clock(clock), .in1(R7710));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7761 (.out1(R7762), .clock(clock), .in1(R7761));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7808 (.out1(R7809), .clock(clock), .in1(R7808));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7861 (.out1(R7862), .clock(clock), .in1(_1029));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7862 (.out1(R7863), .clock(clock), .in1(_1019));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7863 (.out1(R7864), .clock(clock), .in1(_1013));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7864 (.out1(R7865), .clock(clock), .in1(_1001));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7865 (.out1(R7866), .clock(clock), .in1(_995));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7866 (.out1(R7867), .clock(clock), .in1(_985));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7867 (.out1(R7868), .clock(clock), .in1(_1036));
  SRAM op1095 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1037),.ADR(R7868));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1036 (.out1(_978), .in1(R7711));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1037 (.out1(_979), .in1(_978), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1088 (.out1(_1030), .in1(c104_bitmap_2639_D), .in2(R7862));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1078 (.out1(_1020), .in1(c104_bitmap_2639_D), .in2(R7863));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1072 (.out1(_1014), .in1(c104_bitmap_2639_D), .in2(R7864));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1060 (.out1(_1002), .in1(c104_bitmap_2639_D), .in2(R7865));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1054 (.out1(_996), .in1(c104_bitmap_2639_D), .in2(R7866));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1044 (.out1(_986), .in1(c104_bitmap_2639_D), .in2(R7867));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2831 (.out1(R2832), .clock(clock), .in1(R2831));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3037 (.out1(R3038), .clock(clock), .in1(R3037));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3239 (.out1(R3240), .clock(clock), .in1(R3239));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3486 (.out1(R3487), .clock(clock), .in1(R3486));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3678 (.out1(R3679), .clock(clock), .in1(R3678));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3866 (.out1(R3867), .clock(clock), .in1(R3866));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4099 (.out1(R4100), .clock(clock), .in1(R4099));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4277 (.out1(R4278), .clock(clock), .in1(R4277));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4451 (.out1(R4452), .clock(clock), .in1(R4451));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4670 (.out1(R4671), .clock(clock), .in1(R4670));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4834 (.out1(R4835), .clock(clock), .in1(R4834));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4994 (.out1(R4995), .clock(clock), .in1(R4994));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5199 (.out1(R5200), .clock(clock), .in1(R5199));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5349 (.out1(R5350), .clock(clock), .in1(R5349));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5495 (.out1(R5496), .clock(clock), .in1(R5495));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5686 (.out1(R5687), .clock(clock), .in1(R5686));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5822 (.out1(R5823), .clock(clock), .in1(R5822));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5954 (.out1(R5955), .clock(clock), .in1(R5954));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6130 (.out1(R6131), .clock(clock), .in1(R6130));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6251 (.out1(R6252), .clock(clock), .in1(R6251));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6368 (.out1(R6369), .clock(clock), .in1(R6368));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6531 (.out1(R6532), .clock(clock), .in1(R6531));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6638 (.out1(R6639), .clock(clock), .in1(R6638));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6741 (.out1(R6742), .clock(clock), .in1(R6741));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6889 (.out1(R6890), .clock(clock), .in1(R6889));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6982 (.out1(R6983), .clock(clock), .in1(R6982));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7071 (.out1(R7072), .clock(clock), .in1(R7071));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7205 (.out1(R7206), .clock(clock), .in1(R7205));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7284 (.out1(R7285), .clock(clock), .in1(R7284));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7359 (.out1(R7360), .clock(clock), .in1(R7359));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7479 (.out1(R7480), .clock(clock), .in1(R7479));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7544 (.out1(R7545), .clock(clock), .in1(R7544));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7605 (.out1(R7606), .clock(clock), .in1(R7605));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7711 (.out1(R7712), .clock(clock), .in1(R7711));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7762 (.out1(R7763), .clock(clock), .in1(R7762));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7809 (.out1(R7810), .clock(clock), .in1(R7809));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7868 (.out1(R7869), .clock(clock), .in1(_1037));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7869 (.out1(R7870), .clock(clock), .in1(_979));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7870 (.out1(R7871), .clock(clock), .in1(_1030));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7871 (.out1(R7872), .clock(clock), .in1(_1020));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7872 (.out1(R7873), .clock(clock), .in1(_1014));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7873 (.out1(R7874), .clock(clock), .in1(_1002));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7874 (.out1(R7875), .clock(clock), .in1(_996));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7875 (.out1(R7876), .clock(clock), .in1(_986));
  SRAM op1089 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1031),.ADR(R7871));
  SRAM op1079 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1021),.ADR(R7872));
  SRAM op1073 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1015),.ADR(R7873));
  SRAM op1061 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1003),.ADR(R7874));
  SRAM op1055 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_997),.ADR(R7875));
  SRAM op1045 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_987),.ADR(R7876));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1096 (.out1(_1038), .in1(7 'd 64), .in2(R7763));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1038 (.out1(_980), .in1(c104_bitmap_2639_D), .in2(R7870));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1097 (.out1(_1039), .in1(R7869), .in2(_1038));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1090 (.out1(_1032), .in1(7 'd 64), .in2(R7763));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1080 (.out1(_1022), .in1(7 'd 64), .in2(R7763));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1062 (.out1(_1004), .in1(7 'd 64), .in2(R7763));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2832 (.out1(R2833), .clock(clock), .in1(R2832));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3038 (.out1(R3039), .clock(clock), .in1(R3038));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3240 (.out1(R3241), .clock(clock), .in1(R3240));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3487 (.out1(R3488), .clock(clock), .in1(R3487));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3679 (.out1(R3680), .clock(clock), .in1(R3679));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3867 (.out1(R3868), .clock(clock), .in1(R3867));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4100 (.out1(R4101), .clock(clock), .in1(R4100));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4278 (.out1(R4279), .clock(clock), .in1(R4278));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4452 (.out1(R4453), .clock(clock), .in1(R4452));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4671 (.out1(R4672), .clock(clock), .in1(R4671));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4835 (.out1(R4836), .clock(clock), .in1(R4835));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4995 (.out1(R4996), .clock(clock), .in1(R4995));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5200 (.out1(R5201), .clock(clock), .in1(R5200));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5350 (.out1(R5351), .clock(clock), .in1(R5350));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5496 (.out1(R5497), .clock(clock), .in1(R5496));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5687 (.out1(R5688), .clock(clock), .in1(R5687));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5823 (.out1(R5824), .clock(clock), .in1(R5823));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5955 (.out1(R5956), .clock(clock), .in1(R5955));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6131 (.out1(R6132), .clock(clock), .in1(R6131));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6252 (.out1(R6253), .clock(clock), .in1(R6252));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6369 (.out1(R6370), .clock(clock), .in1(R6369));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6532 (.out1(R6533), .clock(clock), .in1(R6532));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6639 (.out1(R6640), .clock(clock), .in1(R6639));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6742 (.out1(R6743), .clock(clock), .in1(R6742));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6890 (.out1(R6891), .clock(clock), .in1(R6890));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6983 (.out1(R6984), .clock(clock), .in1(R6983));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7072 (.out1(R7073), .clock(clock), .in1(R7072));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7206 (.out1(R7207), .clock(clock), .in1(R7206));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7285 (.out1(R7286), .clock(clock), .in1(R7285));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7360 (.out1(R7361), .clock(clock), .in1(R7360));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7480 (.out1(R7481), .clock(clock), .in1(R7480));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7545 (.out1(R7546), .clock(clock), .in1(R7545));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7606 (.out1(R7607), .clock(clock), .in1(R7606));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7712 (.out1(R7713), .clock(clock), .in1(R7712));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7763 (.out1(R7764), .clock(clock), .in1(R7763));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7810 (.out1(R7811), .clock(clock), .in1(R7810));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7876 (.out1(R7877), .clock(clock), .in1(_1031));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7877 (.out1(R7878), .clock(clock), .in1(_1021));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7878 (.out1(R7879), .clock(clock), .in1(_1015));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7879 (.out1(R7880), .clock(clock), .in1(_1003));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7880 (.out1(R7881), .clock(clock), .in1(_997));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7881 (.out1(R7882), .clock(clock), .in1(_987));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7882 (.out1(R7883), .clock(clock), .in1(_980));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7883 (.out1(R7884), .clock(clock), .in1(_1039));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7884 (.out1(R7885), .clock(clock), .in1(_1032));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7885 (.out1(R7886), .clock(clock), .in1(_1022));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7886 (.out1(R7887), .clock(clock), .in1(_1004));
  SRAM op1039 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_981),.ADR(R7883));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1098 (.out1(_1040), .in1(R7884), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1091 (.out1(_1033), .in1(R7877), .in2(R7885));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1081 (.out1(_1023), .in1(R7878), .in2(R7886));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1074 (.out1(_1016), .in1(7 'd 64), .in2(R7764));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1063 (.out1(_1005), .in1(R7880), .in2(R7887));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1056 (.out1(_998), .in1(7 'd 64), .in2(R7764));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1046 (.out1(_988), .in1(7 'd 64), .in2(R7764));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1099 (.out1(_1041), .in1(_1040), .in2(63 'd 6148914691236517205));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1100 (.out1(_1042), .in1(_1033), .in2(_1041));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1082 (.out1(_1024), .in1(_1023), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1075 (.out1(_1017), .in1(R7879), .in2(_1016));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1064 (.out1(_1006), .in1(_1005), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1057 (.out1(_999), .in1(R7881), .in2(_998));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1047 (.out1(_989), .in1(R7882), .in2(_988));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1040 (.out1(_982), .in1(7 'd 64), .in2(R7764));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2833 (.out1(R2834), .clock(clock), .in1(R2833));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3039 (.out1(R3040), .clock(clock), .in1(R3039));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3241 (.out1(R3242), .clock(clock), .in1(R3241));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3488 (.out1(R3489), .clock(clock), .in1(R3488));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3680 (.out1(R3681), .clock(clock), .in1(R3680));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3868 (.out1(R3869), .clock(clock), .in1(R3868));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4101 (.out1(R4102), .clock(clock), .in1(R4101));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4279 (.out1(R4280), .clock(clock), .in1(R4279));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4453 (.out1(R4454), .clock(clock), .in1(R4453));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4672 (.out1(R4673), .clock(clock), .in1(R4672));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4836 (.out1(R4837), .clock(clock), .in1(R4836));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4996 (.out1(R4997), .clock(clock), .in1(R4996));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5201 (.out1(R5202), .clock(clock), .in1(R5201));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5351 (.out1(R5352), .clock(clock), .in1(R5351));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5497 (.out1(R5498), .clock(clock), .in1(R5497));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5688 (.out1(R5689), .clock(clock), .in1(R5688));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5824 (.out1(R5825), .clock(clock), .in1(R5824));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5956 (.out1(R5957), .clock(clock), .in1(R5956));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6132 (.out1(R6133), .clock(clock), .in1(R6132));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6253 (.out1(R6254), .clock(clock), .in1(R6253));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6370 (.out1(R6371), .clock(clock), .in1(R6370));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6533 (.out1(R6534), .clock(clock), .in1(R6533));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6640 (.out1(R6641), .clock(clock), .in1(R6640));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6743 (.out1(R6744), .clock(clock), .in1(R6743));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6891 (.out1(R6892), .clock(clock), .in1(R6891));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6984 (.out1(R6985), .clock(clock), .in1(R6984));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7073 (.out1(R7074), .clock(clock), .in1(R7073));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7207 (.out1(R7208), .clock(clock), .in1(R7207));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7286 (.out1(R7287), .clock(clock), .in1(R7286));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7361 (.out1(R7362), .clock(clock), .in1(R7361));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7481 (.out1(R7482), .clock(clock), .in1(R7481));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7546 (.out1(R7547), .clock(clock), .in1(R7546));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7607 (.out1(R7608), .clock(clock), .in1(R7607));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7713 (.out1(R7714), .clock(clock), .in1(R7713));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7764 (.out1(R7765), .clock(clock), .in1(R7764));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7811 (.out1(R7812), .clock(clock), .in1(R7811));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7887 (.out1(R7888), .clock(clock), .in1(_981));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7888 (.out1(R7889), .clock(clock), .in1(_1042));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7889 (.out1(R7890), .clock(clock), .in1(_1024));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7890 (.out1(R7891), .clock(clock), .in1(_1017));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7891 (.out1(R7892), .clock(clock), .in1(_1006));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7892 (.out1(R7893), .clock(clock), .in1(_999));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7893 (.out1(R7894), .clock(clock), .in1(_989));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7894 (.out1(R7895), .clock(clock), .in1(_982));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1032 (.out1(_974), .in1(R7714));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1083 (.out1(_1025), .in1(R7890), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1101 (.out1(_1043), .in1(R7889), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1084 (.out1(_1026), .in1(R7891), .in2(_1025));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1065 (.out1(_1007), .in1(R7892), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1048 (.out1(_990), .in1(R7894), .in2(1 'd 1));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1066 (.out1(_1008), .in1(R7893), .in2(_1007));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1041 (.out1(_983), .in1(R7888), .in2(R7895));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1033 (.out1(_975), .in1(_974), .in2(2 'd 2));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1102 (.out1(_1044), .in1(_1043), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1085 (.out1(_1027), .in1(_1026), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1049 (.out1(_991), .in1(_990), .in2(63 'd 6148914691236517205));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1103 (.out1(_1045), .in1(_1027), .in2(_1044));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1067 (.out1(_1009), .in1(_1008), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1050 (.out1(_992), .in1(_983), .in2(_991));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2834 (.out1(R2835), .clock(clock), .in1(R2834));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3040 (.out1(R3041), .clock(clock), .in1(R3040));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3242 (.out1(R3243), .clock(clock), .in1(R3242));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3489 (.out1(R3490), .clock(clock), .in1(R3489));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3681 (.out1(R3682), .clock(clock), .in1(R3681));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3869 (.out1(R3870), .clock(clock), .in1(R3869));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4102 (.out1(R4103), .clock(clock), .in1(R4102));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4280 (.out1(R4281), .clock(clock), .in1(R4280));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4454 (.out1(R4455), .clock(clock), .in1(R4454));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4673 (.out1(R4674), .clock(clock), .in1(R4673));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4837 (.out1(R4838), .clock(clock), .in1(R4837));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4997 (.out1(R4998), .clock(clock), .in1(R4997));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5202 (.out1(R5203), .clock(clock), .in1(R5202));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5352 (.out1(R5353), .clock(clock), .in1(R5352));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5498 (.out1(R5499), .clock(clock), .in1(R5498));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5689 (.out1(R5690), .clock(clock), .in1(R5689));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5825 (.out1(R5826), .clock(clock), .in1(R5825));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5957 (.out1(R5958), .clock(clock), .in1(R5957));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6133 (.out1(R6134), .clock(clock), .in1(R6133));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6254 (.out1(R6255), .clock(clock), .in1(R6254));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6371 (.out1(R6372), .clock(clock), .in1(R6371));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6534 (.out1(R6535), .clock(clock), .in1(R6534));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6641 (.out1(R6642), .clock(clock), .in1(R6641));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6744 (.out1(R6745), .clock(clock), .in1(R6744));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6892 (.out1(R6893), .clock(clock), .in1(R6892));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6985 (.out1(R6986), .clock(clock), .in1(R6985));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7074 (.out1(R7075), .clock(clock), .in1(R7074));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7208 (.out1(R7209), .clock(clock), .in1(R7208));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7287 (.out1(R7288), .clock(clock), .in1(R7287));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7362 (.out1(R7363), .clock(clock), .in1(R7362));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7482 (.out1(R7483), .clock(clock), .in1(R7482));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7547 (.out1(R7548), .clock(clock), .in1(R7547));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7608 (.out1(R7609), .clock(clock), .in1(R7608));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7714 (.out1(R7715), .clock(clock), .in1(R7714));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7765 (.out1(R7766), .clock(clock), .in1(R7765));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7812 (.out1(R7813), .clock(clock), .in1(R7812));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7895 (.out1(R7896), .clock(clock), .in1(_975));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7896 (.out1(R7897), .clock(clock), .in1(_1045));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7897 (.out1(R7898), .clock(clock), .in1(_1009));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7898 (.out1(R7899), .clock(clock), .in1(_992));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1068 (.out1(_1010), .in1(R7898), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1051 (.out1(_993), .in1(R7899), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op1104 (.out1(_1046), .in1(R7897), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1069 (.out1(_1011), .in1(_993), .in2(_1010));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1034 (.out1(_976), .in1(c104_popcnt_2644_D), .in2(R7896));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1105 (.out1(_1047), .in1(_1011), .in2(_1046));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op1106 (.out1(_1048), .in1(_1047), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2835 (.out1(R2836), .clock(clock), .in1(R2835));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3041 (.out1(R3042), .clock(clock), .in1(R3041));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3243 (.out1(R3244), .clock(clock), .in1(R3243));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3490 (.out1(R3491), .clock(clock), .in1(R3490));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3682 (.out1(R3683), .clock(clock), .in1(R3682));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3870 (.out1(R3871), .clock(clock), .in1(R3870));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4103 (.out1(R4104), .clock(clock), .in1(R4103));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4281 (.out1(R4282), .clock(clock), .in1(R4281));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4455 (.out1(R4456), .clock(clock), .in1(R4455));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4674 (.out1(R4675), .clock(clock), .in1(R4674));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4838 (.out1(R4839), .clock(clock), .in1(R4838));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4998 (.out1(R4999), .clock(clock), .in1(R4998));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5203 (.out1(R5204), .clock(clock), .in1(R5203));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5353 (.out1(R5354), .clock(clock), .in1(R5353));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5499 (.out1(R5500), .clock(clock), .in1(R5499));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5690 (.out1(R5691), .clock(clock), .in1(R5690));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5826 (.out1(R5827), .clock(clock), .in1(R5826));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5958 (.out1(R5959), .clock(clock), .in1(R5958));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6134 (.out1(R6135), .clock(clock), .in1(R6134));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6255 (.out1(R6256), .clock(clock), .in1(R6255));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6372 (.out1(R6373), .clock(clock), .in1(R6372));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6535 (.out1(R6536), .clock(clock), .in1(R6535));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6642 (.out1(R6643), .clock(clock), .in1(R6642));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6745 (.out1(R6746), .clock(clock), .in1(R6745));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6893 (.out1(R6894), .clock(clock), .in1(R6893));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6986 (.out1(R6987), .clock(clock), .in1(R6986));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7075 (.out1(R7076), .clock(clock), .in1(R7075));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7209 (.out1(R7210), .clock(clock), .in1(R7209));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7288 (.out1(R7289), .clock(clock), .in1(R7288));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7363 (.out1(R7364), .clock(clock), .in1(R7363));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7483 (.out1(R7484), .clock(clock), .in1(R7483));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7548 (.out1(R7549), .clock(clock), .in1(R7548));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7609 (.out1(R7610), .clock(clock), .in1(R7609));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7715 (.out1(R7716), .clock(clock), .in1(R7715));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7766 (.out1(R7767), .clock(clock), .in1(R7766));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7813 (.out1(R7814), .clock(clock), .in1(R7813));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7899 (.out1(R7900), .clock(clock), .in1(_976));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7900 (.out1(R7901), .clock(clock), .in1(_1048));
  SRAM op1035 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_977),.ADR(R7900));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op1107 (.out1(_1049), .in1(R7901), .in2(57 'd 72340172838076673));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2836 (.out1(R2837), .clock(clock), .in1(R2836));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3042 (.out1(R3043), .clock(clock), .in1(R3042));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3244 (.out1(R3245), .clock(clock), .in1(R3244));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3491 (.out1(R3492), .clock(clock), .in1(R3491));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3683 (.out1(R3684), .clock(clock), .in1(R3683));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3871 (.out1(R3872), .clock(clock), .in1(R3871));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4104 (.out1(R4105), .clock(clock), .in1(R4104));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4282 (.out1(R4283), .clock(clock), .in1(R4282));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4456 (.out1(R4457), .clock(clock), .in1(R4456));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4675 (.out1(R4676), .clock(clock), .in1(R4675));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4839 (.out1(R4840), .clock(clock), .in1(R4839));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4999 (.out1(R5000), .clock(clock), .in1(R4999));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5204 (.out1(R5205), .clock(clock), .in1(R5204));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5354 (.out1(R5355), .clock(clock), .in1(R5354));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5500 (.out1(R5501), .clock(clock), .in1(R5500));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5691 (.out1(R5692), .clock(clock), .in1(R5691));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5827 (.out1(R5828), .clock(clock), .in1(R5827));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5959 (.out1(R5960), .clock(clock), .in1(R5959));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6135 (.out1(R6136), .clock(clock), .in1(R6135));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6256 (.out1(R6257), .clock(clock), .in1(R6256));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6373 (.out1(R6374), .clock(clock), .in1(R6373));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6536 (.out1(R6537), .clock(clock), .in1(R6536));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6643 (.out1(R6644), .clock(clock), .in1(R6643));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6746 (.out1(R6747), .clock(clock), .in1(R6746));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6894 (.out1(R6895), .clock(clock), .in1(R6894));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6987 (.out1(R6988), .clock(clock), .in1(R6987));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7076 (.out1(R7077), .clock(clock), .in1(R7076));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7210 (.out1(R7211), .clock(clock), .in1(R7210));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7289 (.out1(R7290), .clock(clock), .in1(R7289));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7364 (.out1(R7365), .clock(clock), .in1(R7364));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7484 (.out1(R7485), .clock(clock), .in1(R7484));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7549 (.out1(R7550), .clock(clock), .in1(R7549));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7610 (.out1(R7611), .clock(clock), .in1(R7610));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7716 (.out1(R7717), .clock(clock), .in1(R7716));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7767 (.out1(R7768), .clock(clock), .in1(R7767));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7814 (.out1(R7815), .clock(clock), .in1(R7814));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7901 (.out1(R7902), .clock(clock), .in1(_977));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7902 (.out1(R7903), .clock(clock), .in1(_1049));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op1108 (.out1(_1050), .in1(R7903), .in2(6 'd 56));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1109 (.out1(_1051), .in1(_1050));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1110 (.out1(ck_idx_2645), .in1(R7902), .in2(_1051));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2837 (.out1(R2838), .clock(clock), .in1(R2837));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3043 (.out1(R3044), .clock(clock), .in1(R3043));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3245 (.out1(R3246), .clock(clock), .in1(R3245));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3492 (.out1(R3493), .clock(clock), .in1(R3492));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3684 (.out1(R3685), .clock(clock), .in1(R3684));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3872 (.out1(R3873), .clock(clock), .in1(R3872));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4105 (.out1(R4106), .clock(clock), .in1(R4105));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4283 (.out1(R4284), .clock(clock), .in1(R4283));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4457 (.out1(R4458), .clock(clock), .in1(R4457));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4676 (.out1(R4677), .clock(clock), .in1(R4676));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4840 (.out1(R4841), .clock(clock), .in1(R4840));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5000 (.out1(R5001), .clock(clock), .in1(R5000));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5205 (.out1(R5206), .clock(clock), .in1(R5205));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5355 (.out1(R5356), .clock(clock), .in1(R5355));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5501 (.out1(R5502), .clock(clock), .in1(R5501));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5692 (.out1(R5693), .clock(clock), .in1(R5692));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5828 (.out1(R5829), .clock(clock), .in1(R5828));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5960 (.out1(R5961), .clock(clock), .in1(R5960));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6136 (.out1(R6137), .clock(clock), .in1(R6136));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6257 (.out1(R6258), .clock(clock), .in1(R6257));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6374 (.out1(R6375), .clock(clock), .in1(R6374));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6537 (.out1(R6538), .clock(clock), .in1(R6537));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6644 (.out1(R6645), .clock(clock), .in1(R6644));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6747 (.out1(R6748), .clock(clock), .in1(R6747));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6895 (.out1(R6896), .clock(clock), .in1(R6895));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6988 (.out1(R6989), .clock(clock), .in1(R6988));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7077 (.out1(R7078), .clock(clock), .in1(R7077));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7211 (.out1(R7212), .clock(clock), .in1(R7211));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7290 (.out1(R7291), .clock(clock), .in1(R7290));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7365 (.out1(R7366), .clock(clock), .in1(R7365));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7485 (.out1(R7486), .clock(clock), .in1(R7485));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7550 (.out1(R7551), .clock(clock), .in1(R7550));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7611 (.out1(R7612), .clock(clock), .in1(R7611));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7717 (.out1(R7718), .clock(clock), .in1(R7717));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7768 (.out1(R7769), .clock(clock), .in1(R7768));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7815 (.out1(R7816), .clock(clock), .in1(R7815));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7903 (.out1(R7904), .clock(clock), .in1(ck_idx_2645));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(4), .BITSIZE_out1(32), .PRECISION(32)) op1111 (.out1(_1052), .in1(R7904), .in2(4 'd 8));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(5), .BITSIZE_out1(64), .PRECISION(64)) op1112 (.out1(_1053), .in1(ip2_2595_D), .in2(5 'd 16));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2838 (.out1(R2839), .clock(clock), .in1(R2838));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3044 (.out1(R3045), .clock(clock), .in1(R3044));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3246 (.out1(R3247), .clock(clock), .in1(R3246));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3493 (.out1(R3494), .clock(clock), .in1(R3493));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3685 (.out1(R3686), .clock(clock), .in1(R3685));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3873 (.out1(R3874), .clock(clock), .in1(R3873));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4106 (.out1(R4107), .clock(clock), .in1(R4106));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4284 (.out1(R4285), .clock(clock), .in1(R4284));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4458 (.out1(R4459), .clock(clock), .in1(R4458));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4677 (.out1(R4678), .clock(clock), .in1(R4677));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4841 (.out1(R4842), .clock(clock), .in1(R4841));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5001 (.out1(R5002), .clock(clock), .in1(R5001));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5206 (.out1(R5207), .clock(clock), .in1(R5206));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5356 (.out1(R5357), .clock(clock), .in1(R5356));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5502 (.out1(R5503), .clock(clock), .in1(R5502));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5693 (.out1(R5694), .clock(clock), .in1(R5693));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5829 (.out1(R5830), .clock(clock), .in1(R5829));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5961 (.out1(R5962), .clock(clock), .in1(R5961));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6137 (.out1(R6138), .clock(clock), .in1(R6137));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6258 (.out1(R6259), .clock(clock), .in1(R6258));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6375 (.out1(R6376), .clock(clock), .in1(R6375));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6538 (.out1(R6539), .clock(clock), .in1(R6538));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6645 (.out1(R6646), .clock(clock), .in1(R6645));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6748 (.out1(R6749), .clock(clock), .in1(R6748));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6896 (.out1(R6897), .clock(clock), .in1(R6896));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6989 (.out1(R6990), .clock(clock), .in1(R6989));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7078 (.out1(R7079), .clock(clock), .in1(R7078));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7212 (.out1(R7213), .clock(clock), .in1(R7212));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7291 (.out1(R7292), .clock(clock), .in1(R7291));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7366 (.out1(R7367), .clock(clock), .in1(R7366));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7486 (.out1(R7487), .clock(clock), .in1(R7486));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7551 (.out1(R7552), .clock(clock), .in1(R7551));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7612 (.out1(R7613), .clock(clock), .in1(R7612));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7718 (.out1(R7719), .clock(clock), .in1(R7718));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7769 (.out1(R7770), .clock(clock), .in1(R7769));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7816 (.out1(R7817), .clock(clock), .in1(R7816));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7904 (.out1(R7905), .clock(clock), .in1(_1052));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7905 (.out1(R7906), .clock(clock), .in1(_1053));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1113 (.out1(_1054), .in1(R7906));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(8), .BITSIZE_out1(32)) op1114 (.out1(_1055), .in1(_1054), .in2(8 'd 255));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1115 (.out1(idx_sail_2646), .in1(R7905), .in2(_1055));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(3), .BITSIZE_out1(32), .PRECISION(32)) op1116 (.out1(idx_2647), .in1(idx_sail_2646), .in2(3 'd 6));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2839 (.out1(R2840), .clock(clock), .in1(R2839));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3045 (.out1(R3046), .clock(clock), .in1(R3045));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3247 (.out1(R3248), .clock(clock), .in1(R3247));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3494 (.out1(R3495), .clock(clock), .in1(R3494));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3686 (.out1(R3687), .clock(clock), .in1(R3686));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3874 (.out1(R3875), .clock(clock), .in1(R3874));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4107 (.out1(R4108), .clock(clock), .in1(R4107));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4285 (.out1(R4286), .clock(clock), .in1(R4285));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4459 (.out1(R4460), .clock(clock), .in1(R4459));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4678 (.out1(R4679), .clock(clock), .in1(R4678));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4842 (.out1(R4843), .clock(clock), .in1(R4842));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5002 (.out1(R5003), .clock(clock), .in1(R5002));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5207 (.out1(R5208), .clock(clock), .in1(R5207));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5357 (.out1(R5358), .clock(clock), .in1(R5357));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5503 (.out1(R5504), .clock(clock), .in1(R5503));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5694 (.out1(R5695), .clock(clock), .in1(R5694));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5830 (.out1(R5831), .clock(clock), .in1(R5830));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5962 (.out1(R5963), .clock(clock), .in1(R5962));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6138 (.out1(R6139), .clock(clock), .in1(R6138));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6259 (.out1(R6260), .clock(clock), .in1(R6259));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6376 (.out1(R6377), .clock(clock), .in1(R6376));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6539 (.out1(R6540), .clock(clock), .in1(R6539));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6646 (.out1(R6647), .clock(clock), .in1(R6646));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6749 (.out1(R6750), .clock(clock), .in1(R6749));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6897 (.out1(R6898), .clock(clock), .in1(R6897));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6990 (.out1(R6991), .clock(clock), .in1(R6990));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7079 (.out1(R7080), .clock(clock), .in1(R7079));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7213 (.out1(R7214), .clock(clock), .in1(R7213));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7292 (.out1(R7293), .clock(clock), .in1(R7292));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7367 (.out1(R7368), .clock(clock), .in1(R7367));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7487 (.out1(R7488), .clock(clock), .in1(R7487));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7552 (.out1(R7553), .clock(clock), .in1(R7552));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7613 (.out1(R7614), .clock(clock), .in1(R7613));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7719 (.out1(R7720), .clock(clock), .in1(R7719));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7770 (.out1(R7771), .clock(clock), .in1(R7770));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7817 (.out1(R7818), .clock(clock), .in1(R7817));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7906 (.out1(R7907), .clock(clock), .in1(idx_sail_2646));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7909 (.out1(R7910), .clock(clock), .in1(idx_2647));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1118 (.out1(_1056), .in1(R7910));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1119 (.out1(_1057), .in1(_1056), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2840 (.out1(R2841), .clock(clock), .in1(R2840));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3046 (.out1(R3047), .clock(clock), .in1(R3046));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3248 (.out1(R3249), .clock(clock), .in1(R3248));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3495 (.out1(R3496), .clock(clock), .in1(R3495));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3687 (.out1(R3688), .clock(clock), .in1(R3687));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3875 (.out1(R3876), .clock(clock), .in1(R3875));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4108 (.out1(R4109), .clock(clock), .in1(R4108));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4286 (.out1(R4287), .clock(clock), .in1(R4286));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4460 (.out1(R4461), .clock(clock), .in1(R4460));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4679 (.out1(R4680), .clock(clock), .in1(R4679));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4843 (.out1(R4844), .clock(clock), .in1(R4843));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5003 (.out1(R5004), .clock(clock), .in1(R5003));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5208 (.out1(R5209), .clock(clock), .in1(R5208));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5358 (.out1(R5359), .clock(clock), .in1(R5358));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5504 (.out1(R5505), .clock(clock), .in1(R5504));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5695 (.out1(R5696), .clock(clock), .in1(R5695));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5831 (.out1(R5832), .clock(clock), .in1(R5831));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5963 (.out1(R5964), .clock(clock), .in1(R5963));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6139 (.out1(R6140), .clock(clock), .in1(R6139));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6260 (.out1(R6261), .clock(clock), .in1(R6260));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6377 (.out1(R6378), .clock(clock), .in1(R6377));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6540 (.out1(R6541), .clock(clock), .in1(R6540));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6647 (.out1(R6648), .clock(clock), .in1(R6647));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6750 (.out1(R6751), .clock(clock), .in1(R6750));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6898 (.out1(R6899), .clock(clock), .in1(R6898));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6991 (.out1(R6992), .clock(clock), .in1(R6991));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7080 (.out1(R7081), .clock(clock), .in1(R7080));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7214 (.out1(R7215), .clock(clock), .in1(R7214));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7293 (.out1(R7294), .clock(clock), .in1(R7293));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7368 (.out1(R7369), .clock(clock), .in1(R7368));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7488 (.out1(R7489), .clock(clock), .in1(R7488));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7553 (.out1(R7554), .clock(clock), .in1(R7553));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7614 (.out1(R7615), .clock(clock), .in1(R7614));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7720 (.out1(R7721), .clock(clock), .in1(R7720));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7771 (.out1(R7772), .clock(clock), .in1(R7771));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7818 (.out1(R7819), .clock(clock), .in1(R7818));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7907 (.out1(R7908), .clock(clock), .in1(R7907));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7910 (.out1(R7911), .clock(clock), .in1(R7910));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7946 (.out1(R7947), .clock(clock), .in1(_1057));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1120 (.out1(_1058), .in1(c112_bitmap_2649_D), .in2(R7947));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2841 (.out1(R2842), .clock(clock), .in1(R2841));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3047 (.out1(R3048), .clock(clock), .in1(R3047));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3249 (.out1(R3250), .clock(clock), .in1(R3249));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3496 (.out1(R3497), .clock(clock), .in1(R3496));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3688 (.out1(R3689), .clock(clock), .in1(R3688));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3876 (.out1(R3877), .clock(clock), .in1(R3876));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4109 (.out1(R4110), .clock(clock), .in1(R4109));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4287 (.out1(R4288), .clock(clock), .in1(R4287));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4461 (.out1(R4462), .clock(clock), .in1(R4461));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4680 (.out1(R4681), .clock(clock), .in1(R4680));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4844 (.out1(R4845), .clock(clock), .in1(R4844));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5004 (.out1(R5005), .clock(clock), .in1(R5004));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5209 (.out1(R5210), .clock(clock), .in1(R5209));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5359 (.out1(R5360), .clock(clock), .in1(R5359));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5505 (.out1(R5506), .clock(clock), .in1(R5505));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5696 (.out1(R5697), .clock(clock), .in1(R5696));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5832 (.out1(R5833), .clock(clock), .in1(R5832));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5964 (.out1(R5965), .clock(clock), .in1(R5964));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6140 (.out1(R6141), .clock(clock), .in1(R6140));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6261 (.out1(R6262), .clock(clock), .in1(R6261));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6378 (.out1(R6379), .clock(clock), .in1(R6378));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6541 (.out1(R6542), .clock(clock), .in1(R6541));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6648 (.out1(R6649), .clock(clock), .in1(R6648));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6751 (.out1(R6752), .clock(clock), .in1(R6751));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6899 (.out1(R6900), .clock(clock), .in1(R6899));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6992 (.out1(R6993), .clock(clock), .in1(R6992));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7081 (.out1(R7082), .clock(clock), .in1(R7081));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7215 (.out1(R7216), .clock(clock), .in1(R7215));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7294 (.out1(R7295), .clock(clock), .in1(R7294));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7369 (.out1(R7370), .clock(clock), .in1(R7369));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7489 (.out1(R7490), .clock(clock), .in1(R7489));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7554 (.out1(R7555), .clock(clock), .in1(R7554));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7615 (.out1(R7616), .clock(clock), .in1(R7615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7721 (.out1(R7722), .clock(clock), .in1(R7721));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7772 (.out1(R7773), .clock(clock), .in1(R7772));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7819 (.out1(R7820), .clock(clock), .in1(R7819));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7908 (.out1(R7909), .clock(clock), .in1(R7908));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7911 (.out1(R7912), .clock(clock), .in1(R7911));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7947 (.out1(R7948), .clock(clock), .in1(_1058));
  SRAM op1121 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1059),.ADR(R7948));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op1117 (.out1(off_2648), .in1(R7909), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1122 (.out1(_1060), .in1(64 'd 9223372036854775808), .in2(off_2648));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2842 (.out1(R2843), .clock(clock), .in1(R2842));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3048 (.out1(R3049), .clock(clock), .in1(R3048));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3250 (.out1(R3251), .clock(clock), .in1(R3250));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3497 (.out1(R3498), .clock(clock), .in1(R3497));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3689 (.out1(R3690), .clock(clock), .in1(R3689));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3877 (.out1(R3878), .clock(clock), .in1(R3877));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4110 (.out1(R4111), .clock(clock), .in1(R4110));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4288 (.out1(R4289), .clock(clock), .in1(R4288));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4462 (.out1(R4463), .clock(clock), .in1(R4462));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4681 (.out1(R4682), .clock(clock), .in1(R4681));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4845 (.out1(R4846), .clock(clock), .in1(R4845));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5005 (.out1(R5006), .clock(clock), .in1(R5005));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5210 (.out1(R5211), .clock(clock), .in1(R5210));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5360 (.out1(R5361), .clock(clock), .in1(R5360));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5506 (.out1(R5507), .clock(clock), .in1(R5506));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5697 (.out1(R5698), .clock(clock), .in1(R5697));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5833 (.out1(R5834), .clock(clock), .in1(R5833));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5965 (.out1(R5966), .clock(clock), .in1(R5965));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6141 (.out1(R6142), .clock(clock), .in1(R6141));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6262 (.out1(R6263), .clock(clock), .in1(R6262));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6379 (.out1(R6380), .clock(clock), .in1(R6379));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6542 (.out1(R6543), .clock(clock), .in1(R6542));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6649 (.out1(R6650), .clock(clock), .in1(R6649));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6752 (.out1(R6753), .clock(clock), .in1(R6752));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6900 (.out1(R6901), .clock(clock), .in1(R6900));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6993 (.out1(R6994), .clock(clock), .in1(R6993));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7082 (.out1(R7083), .clock(clock), .in1(R7082));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7216 (.out1(R7217), .clock(clock), .in1(R7216));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7295 (.out1(R7296), .clock(clock), .in1(R7295));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7370 (.out1(R7371), .clock(clock), .in1(R7370));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7490 (.out1(R7491), .clock(clock), .in1(R7490));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7555 (.out1(R7556), .clock(clock), .in1(R7555));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7616 (.out1(R7617), .clock(clock), .in1(R7616));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7722 (.out1(R7723), .clock(clock), .in1(R7722));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7773 (.out1(R7774), .clock(clock), .in1(R7773));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7820 (.out1(R7821), .clock(clock), .in1(R7820));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7912 (.out1(R7913), .clock(clock), .in1(R7912));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7948 (.out1(R7949), .clock(clock), .in1(_1059));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7949 (.out1(R7950), .clock(clock), .in1(off_2648));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7982 (.out1(R7983), .clock(clock), .in1(_1060));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1123 (.out1(_1061), .in1(R7949), .in2(R7983));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op1124 (.out1(ifout1124), .in1(_1061), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1185 (.out1(_1122), .in1(R7913));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1186 (.out1(_1123), .in1(_1122), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2843 (.out1(R2844), .clock(clock), .in1(R2843));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3049 (.out1(R3050), .clock(clock), .in1(R3049));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3251 (.out1(R3252), .clock(clock), .in1(R3251));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3498 (.out1(R3499), .clock(clock), .in1(R3498));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3690 (.out1(R3691), .clock(clock), .in1(R3690));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3878 (.out1(R3879), .clock(clock), .in1(R3878));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4111 (.out1(R4112), .clock(clock), .in1(R4111));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4289 (.out1(R4290), .clock(clock), .in1(R4289));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4463 (.out1(R4464), .clock(clock), .in1(R4463));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4682 (.out1(R4683), .clock(clock), .in1(R4682));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4846 (.out1(R4847), .clock(clock), .in1(R4846));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5006 (.out1(R5007), .clock(clock), .in1(R5006));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5211 (.out1(R5212), .clock(clock), .in1(R5211));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5361 (.out1(R5362), .clock(clock), .in1(R5361));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5507 (.out1(R5508), .clock(clock), .in1(R5507));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5698 (.out1(R5699), .clock(clock), .in1(R5698));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5834 (.out1(R5835), .clock(clock), .in1(R5834));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5966 (.out1(R5967), .clock(clock), .in1(R5966));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6142 (.out1(R6143), .clock(clock), .in1(R6142));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6263 (.out1(R6264), .clock(clock), .in1(R6263));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6380 (.out1(R6381), .clock(clock), .in1(R6380));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6543 (.out1(R6544), .clock(clock), .in1(R6543));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6650 (.out1(R6651), .clock(clock), .in1(R6650));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6753 (.out1(R6754), .clock(clock), .in1(R6753));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6901 (.out1(R6902), .clock(clock), .in1(R6901));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6994 (.out1(R6995), .clock(clock), .in1(R6994));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7083 (.out1(R7084), .clock(clock), .in1(R7083));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7217 (.out1(R7218), .clock(clock), .in1(R7217));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7296 (.out1(R7297), .clock(clock), .in1(R7296));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7371 (.out1(R7372), .clock(clock), .in1(R7371));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7491 (.out1(R7492), .clock(clock), .in1(R7491));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7556 (.out1(R7557), .clock(clock), .in1(R7556));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7617 (.out1(R7618), .clock(clock), .in1(R7617));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7723 (.out1(R7724), .clock(clock), .in1(R7723));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7774 (.out1(R7775), .clock(clock), .in1(R7774));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7821 (.out1(R7822), .clock(clock), .in1(R7821));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7913 (.out1(R7914), .clock(clock), .in1(R7913));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7950 (.out1(R7951), .clock(clock), .in1(R7950));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7983 (.out1(R7984), .clock(clock), .in1(ifout1124));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8022 (.out1(R8023), .clock(clock), .in1(_1123));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1179 (.out1(_1116), .in1(R7914));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1169 (.out1(_1106), .in1(R7914));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1163 (.out1(_1100), .in1(R7914));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1151 (.out1(_1088), .in1(R7914));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1145 (.out1(_1082), .in1(R7914));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1135 (.out1(_1072), .in1(R7914));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1180 (.out1(_1117), .in1(_1116), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1170 (.out1(_1107), .in1(_1106), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1164 (.out1(_1101), .in1(_1100), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1152 (.out1(_1089), .in1(_1088), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1146 (.out1(_1083), .in1(_1082), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1136 (.out1(_1073), .in1(_1072), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1187 (.out1(_1124), .in1(c112_bitmap_2649_D), .in2(R8023));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2844 (.out1(R2845), .clock(clock), .in1(R2844));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3050 (.out1(R3051), .clock(clock), .in1(R3050));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3252 (.out1(R3253), .clock(clock), .in1(R3252));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3499 (.out1(R3500), .clock(clock), .in1(R3499));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3691 (.out1(R3692), .clock(clock), .in1(R3691));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3879 (.out1(R3880), .clock(clock), .in1(R3879));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4112 (.out1(R4113), .clock(clock), .in1(R4112));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4290 (.out1(R4291), .clock(clock), .in1(R4290));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4464 (.out1(R4465), .clock(clock), .in1(R4464));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4683 (.out1(R4684), .clock(clock), .in1(R4683));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4847 (.out1(R4848), .clock(clock), .in1(R4847));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5007 (.out1(R5008), .clock(clock), .in1(R5007));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5212 (.out1(R5213), .clock(clock), .in1(R5212));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5362 (.out1(R5363), .clock(clock), .in1(R5362));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5508 (.out1(R5509), .clock(clock), .in1(R5508));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5699 (.out1(R5700), .clock(clock), .in1(R5699));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5835 (.out1(R5836), .clock(clock), .in1(R5835));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5967 (.out1(R5968), .clock(clock), .in1(R5967));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6143 (.out1(R6144), .clock(clock), .in1(R6143));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6264 (.out1(R6265), .clock(clock), .in1(R6264));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6381 (.out1(R6382), .clock(clock), .in1(R6381));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6544 (.out1(R6545), .clock(clock), .in1(R6544));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6651 (.out1(R6652), .clock(clock), .in1(R6651));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6754 (.out1(R6755), .clock(clock), .in1(R6754));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6902 (.out1(R6903), .clock(clock), .in1(R6902));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6995 (.out1(R6996), .clock(clock), .in1(R6995));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7084 (.out1(R7085), .clock(clock), .in1(R7084));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7218 (.out1(R7219), .clock(clock), .in1(R7218));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7297 (.out1(R7298), .clock(clock), .in1(R7297));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7372 (.out1(R7373), .clock(clock), .in1(R7372));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7492 (.out1(R7493), .clock(clock), .in1(R7492));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7557 (.out1(R7558), .clock(clock), .in1(R7557));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7618 (.out1(R7619), .clock(clock), .in1(R7618));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7724 (.out1(R7725), .clock(clock), .in1(R7724));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7775 (.out1(R7776), .clock(clock), .in1(R7775));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7822 (.out1(R7823), .clock(clock), .in1(R7822));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7914 (.out1(R7915), .clock(clock), .in1(R7914));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7951 (.out1(R7952), .clock(clock), .in1(R7951));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7984 (.out1(R7985), .clock(clock), .in1(R7984));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8023 (.out1(R8024), .clock(clock), .in1(_1117));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8024 (.out1(R8025), .clock(clock), .in1(_1107));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8025 (.out1(R8026), .clock(clock), .in1(_1101));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8026 (.out1(R8027), .clock(clock), .in1(_1089));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8027 (.out1(R8028), .clock(clock), .in1(_1083));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8028 (.out1(R8029), .clock(clock), .in1(_1073));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8029 (.out1(R8030), .clock(clock), .in1(_1124));
  SRAM op1188 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1125),.ADR(R8030));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1129 (.out1(_1066), .in1(R7915));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1130 (.out1(_1067), .in1(_1066), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1181 (.out1(_1118), .in1(c112_bitmap_2649_D), .in2(R8024));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1171 (.out1(_1108), .in1(c112_bitmap_2649_D), .in2(R8025));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1165 (.out1(_1102), .in1(c112_bitmap_2649_D), .in2(R8026));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1153 (.out1(_1090), .in1(c112_bitmap_2649_D), .in2(R8027));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1147 (.out1(_1084), .in1(c112_bitmap_2649_D), .in2(R8028));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1137 (.out1(_1074), .in1(c112_bitmap_2649_D), .in2(R8029));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2845 (.out1(R2846), .clock(clock), .in1(R2845));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3051 (.out1(R3052), .clock(clock), .in1(R3051));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3253 (.out1(R3254), .clock(clock), .in1(R3253));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3500 (.out1(R3501), .clock(clock), .in1(R3500));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3692 (.out1(R3693), .clock(clock), .in1(R3692));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3880 (.out1(R3881), .clock(clock), .in1(R3880));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4113 (.out1(R4114), .clock(clock), .in1(R4113));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4291 (.out1(R4292), .clock(clock), .in1(R4291));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4465 (.out1(R4466), .clock(clock), .in1(R4465));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4684 (.out1(R4685), .clock(clock), .in1(R4684));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4848 (.out1(R4849), .clock(clock), .in1(R4848));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5008 (.out1(R5009), .clock(clock), .in1(R5008));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5213 (.out1(R5214), .clock(clock), .in1(R5213));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5363 (.out1(R5364), .clock(clock), .in1(R5363));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5509 (.out1(R5510), .clock(clock), .in1(R5509));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5700 (.out1(R5701), .clock(clock), .in1(R5700));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5836 (.out1(R5837), .clock(clock), .in1(R5836));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5968 (.out1(R5969), .clock(clock), .in1(R5968));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6144 (.out1(R6145), .clock(clock), .in1(R6144));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6265 (.out1(R6266), .clock(clock), .in1(R6265));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6382 (.out1(R6383), .clock(clock), .in1(R6382));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6545 (.out1(R6546), .clock(clock), .in1(R6545));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6652 (.out1(R6653), .clock(clock), .in1(R6652));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6755 (.out1(R6756), .clock(clock), .in1(R6755));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6903 (.out1(R6904), .clock(clock), .in1(R6903));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6996 (.out1(R6997), .clock(clock), .in1(R6996));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7085 (.out1(R7086), .clock(clock), .in1(R7085));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7219 (.out1(R7220), .clock(clock), .in1(R7219));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7298 (.out1(R7299), .clock(clock), .in1(R7298));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7373 (.out1(R7374), .clock(clock), .in1(R7373));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7493 (.out1(R7494), .clock(clock), .in1(R7493));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7558 (.out1(R7559), .clock(clock), .in1(R7558));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7619 (.out1(R7620), .clock(clock), .in1(R7619));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7725 (.out1(R7726), .clock(clock), .in1(R7725));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7776 (.out1(R7777), .clock(clock), .in1(R7776));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7823 (.out1(R7824), .clock(clock), .in1(R7823));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7915 (.out1(R7916), .clock(clock), .in1(R7915));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7952 (.out1(R7953), .clock(clock), .in1(R7952));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7985 (.out1(R7986), .clock(clock), .in1(R7985));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8030 (.out1(R8031), .clock(clock), .in1(_1125));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8031 (.out1(R8032), .clock(clock), .in1(_1067));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8032 (.out1(R8033), .clock(clock), .in1(_1118));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8033 (.out1(R8034), .clock(clock), .in1(_1108));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8034 (.out1(R8035), .clock(clock), .in1(_1102));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8035 (.out1(R8036), .clock(clock), .in1(_1090));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8036 (.out1(R8037), .clock(clock), .in1(_1084));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8037 (.out1(R8038), .clock(clock), .in1(_1074));
  SRAM op1182 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1119),.ADR(R8033));
  SRAM op1172 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1109),.ADR(R8034));
  SRAM op1166 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1103),.ADR(R8035));
  SRAM op1154 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1091),.ADR(R8036));
  SRAM op1148 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1085),.ADR(R8037));
  SRAM op1138 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1075),.ADR(R8038));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1189 (.out1(_1126), .in1(7 'd 64), .in2(R7953));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1131 (.out1(_1068), .in1(c112_bitmap_2649_D), .in2(R8032));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1190 (.out1(_1127), .in1(R8031), .in2(_1126));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1183 (.out1(_1120), .in1(7 'd 64), .in2(R7953));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1173 (.out1(_1110), .in1(7 'd 64), .in2(R7953));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1155 (.out1(_1092), .in1(7 'd 64), .in2(R7953));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2846 (.out1(R2847), .clock(clock), .in1(R2846));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3052 (.out1(R3053), .clock(clock), .in1(R3052));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3254 (.out1(R3255), .clock(clock), .in1(R3254));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3501 (.out1(R3502), .clock(clock), .in1(R3501));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3693 (.out1(R3694), .clock(clock), .in1(R3693));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3881 (.out1(R3882), .clock(clock), .in1(R3881));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4114 (.out1(R4115), .clock(clock), .in1(R4114));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4292 (.out1(R4293), .clock(clock), .in1(R4292));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4466 (.out1(R4467), .clock(clock), .in1(R4466));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4685 (.out1(R4686), .clock(clock), .in1(R4685));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4849 (.out1(R4850), .clock(clock), .in1(R4849));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5009 (.out1(R5010), .clock(clock), .in1(R5009));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5214 (.out1(R5215), .clock(clock), .in1(R5214));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5364 (.out1(R5365), .clock(clock), .in1(R5364));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5510 (.out1(R5511), .clock(clock), .in1(R5510));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5701 (.out1(R5702), .clock(clock), .in1(R5701));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5837 (.out1(R5838), .clock(clock), .in1(R5837));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5969 (.out1(R5970), .clock(clock), .in1(R5969));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6145 (.out1(R6146), .clock(clock), .in1(R6145));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6266 (.out1(R6267), .clock(clock), .in1(R6266));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6383 (.out1(R6384), .clock(clock), .in1(R6383));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6546 (.out1(R6547), .clock(clock), .in1(R6546));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6653 (.out1(R6654), .clock(clock), .in1(R6653));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6756 (.out1(R6757), .clock(clock), .in1(R6756));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6904 (.out1(R6905), .clock(clock), .in1(R6904));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6997 (.out1(R6998), .clock(clock), .in1(R6997));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7086 (.out1(R7087), .clock(clock), .in1(R7086));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7220 (.out1(R7221), .clock(clock), .in1(R7220));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7299 (.out1(R7300), .clock(clock), .in1(R7299));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7374 (.out1(R7375), .clock(clock), .in1(R7374));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7494 (.out1(R7495), .clock(clock), .in1(R7494));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7559 (.out1(R7560), .clock(clock), .in1(R7559));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7620 (.out1(R7621), .clock(clock), .in1(R7620));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7726 (.out1(R7727), .clock(clock), .in1(R7726));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7777 (.out1(R7778), .clock(clock), .in1(R7777));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7824 (.out1(R7825), .clock(clock), .in1(R7824));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7916 (.out1(R7917), .clock(clock), .in1(R7916));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7953 (.out1(R7954), .clock(clock), .in1(R7953));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7986 (.out1(R7987), .clock(clock), .in1(R7986));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8038 (.out1(R8039), .clock(clock), .in1(_1119));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8039 (.out1(R8040), .clock(clock), .in1(_1109));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8040 (.out1(R8041), .clock(clock), .in1(_1103));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8041 (.out1(R8042), .clock(clock), .in1(_1091));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8042 (.out1(R8043), .clock(clock), .in1(_1085));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8043 (.out1(R8044), .clock(clock), .in1(_1075));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8044 (.out1(R8045), .clock(clock), .in1(_1068));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8045 (.out1(R8046), .clock(clock), .in1(_1127));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8046 (.out1(R8047), .clock(clock), .in1(_1120));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8047 (.out1(R8048), .clock(clock), .in1(_1110));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8048 (.out1(R8049), .clock(clock), .in1(_1092));
  SRAM op1132 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1069),.ADR(R8045));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1191 (.out1(_1128), .in1(R8046), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1184 (.out1(_1121), .in1(R8039), .in2(R8047));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1174 (.out1(_1111), .in1(R8040), .in2(R8048));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1167 (.out1(_1104), .in1(7 'd 64), .in2(R7954));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1156 (.out1(_1093), .in1(R8042), .in2(R8049));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1149 (.out1(_1086), .in1(7 'd 64), .in2(R7954));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1139 (.out1(_1076), .in1(7 'd 64), .in2(R7954));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1192 (.out1(_1129), .in1(_1128), .in2(63 'd 6148914691236517205));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1193 (.out1(_1130), .in1(_1121), .in2(_1129));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1175 (.out1(_1112), .in1(_1111), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1168 (.out1(_1105), .in1(R8041), .in2(_1104));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1157 (.out1(_1094), .in1(_1093), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1150 (.out1(_1087), .in1(R8043), .in2(_1086));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1140 (.out1(_1077), .in1(R8044), .in2(_1076));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1133 (.out1(_1070), .in1(7 'd 64), .in2(R7954));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2847 (.out1(R2848), .clock(clock), .in1(R2847));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3053 (.out1(R3054), .clock(clock), .in1(R3053));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3255 (.out1(R3256), .clock(clock), .in1(R3255));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3502 (.out1(R3503), .clock(clock), .in1(R3502));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3694 (.out1(R3695), .clock(clock), .in1(R3694));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3882 (.out1(R3883), .clock(clock), .in1(R3882));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4115 (.out1(R4116), .clock(clock), .in1(R4115));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4293 (.out1(R4294), .clock(clock), .in1(R4293));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4467 (.out1(R4468), .clock(clock), .in1(R4467));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4686 (.out1(R4687), .clock(clock), .in1(R4686));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4850 (.out1(R4851), .clock(clock), .in1(R4850));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5010 (.out1(R5011), .clock(clock), .in1(R5010));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5215 (.out1(R5216), .clock(clock), .in1(R5215));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5365 (.out1(R5366), .clock(clock), .in1(R5365));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5511 (.out1(R5512), .clock(clock), .in1(R5511));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5702 (.out1(R5703), .clock(clock), .in1(R5702));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5838 (.out1(R5839), .clock(clock), .in1(R5838));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5970 (.out1(R5971), .clock(clock), .in1(R5970));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6146 (.out1(R6147), .clock(clock), .in1(R6146));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6267 (.out1(R6268), .clock(clock), .in1(R6267));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6384 (.out1(R6385), .clock(clock), .in1(R6384));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6547 (.out1(R6548), .clock(clock), .in1(R6547));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6654 (.out1(R6655), .clock(clock), .in1(R6654));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6757 (.out1(R6758), .clock(clock), .in1(R6757));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6905 (.out1(R6906), .clock(clock), .in1(R6905));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6998 (.out1(R6999), .clock(clock), .in1(R6998));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7087 (.out1(R7088), .clock(clock), .in1(R7087));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7221 (.out1(R7222), .clock(clock), .in1(R7221));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7300 (.out1(R7301), .clock(clock), .in1(R7300));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7375 (.out1(R7376), .clock(clock), .in1(R7375));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7495 (.out1(R7496), .clock(clock), .in1(R7495));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7560 (.out1(R7561), .clock(clock), .in1(R7560));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7621 (.out1(R7622), .clock(clock), .in1(R7621));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7727 (.out1(R7728), .clock(clock), .in1(R7727));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7778 (.out1(R7779), .clock(clock), .in1(R7778));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7825 (.out1(R7826), .clock(clock), .in1(R7825));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7917 (.out1(R7918), .clock(clock), .in1(R7917));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7954 (.out1(R7955), .clock(clock), .in1(R7954));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7987 (.out1(R7988), .clock(clock), .in1(R7987));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8049 (.out1(R8050), .clock(clock), .in1(_1069));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8050 (.out1(R8051), .clock(clock), .in1(_1130));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8051 (.out1(R8052), .clock(clock), .in1(_1112));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8052 (.out1(R8053), .clock(clock), .in1(_1105));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8053 (.out1(R8054), .clock(clock), .in1(_1094));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8054 (.out1(R8055), .clock(clock), .in1(_1087));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8055 (.out1(R8056), .clock(clock), .in1(_1077));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8056 (.out1(R8057), .clock(clock), .in1(_1070));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1125 (.out1(_1062), .in1(R7918));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1176 (.out1(_1113), .in1(R8052), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1194 (.out1(_1131), .in1(R8051), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1177 (.out1(_1114), .in1(R8053), .in2(_1113));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1158 (.out1(_1095), .in1(R8054), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1141 (.out1(_1078), .in1(R8056), .in2(1 'd 1));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1159 (.out1(_1096), .in1(R8055), .in2(_1095));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1134 (.out1(_1071), .in1(R8050), .in2(R8057));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1126 (.out1(_1063), .in1(_1062), .in2(2 'd 2));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1195 (.out1(_1132), .in1(_1131), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1178 (.out1(_1115), .in1(_1114), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1142 (.out1(_1079), .in1(_1078), .in2(63 'd 6148914691236517205));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1196 (.out1(_1133), .in1(_1115), .in2(_1132));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1160 (.out1(_1097), .in1(_1096), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1143 (.out1(_1080), .in1(_1071), .in2(_1079));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2848 (.out1(R2849), .clock(clock), .in1(R2848));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3054 (.out1(R3055), .clock(clock), .in1(R3054));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3256 (.out1(R3257), .clock(clock), .in1(R3256));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3503 (.out1(R3504), .clock(clock), .in1(R3503));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3695 (.out1(R3696), .clock(clock), .in1(R3695));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3883 (.out1(R3884), .clock(clock), .in1(R3883));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4116 (.out1(R4117), .clock(clock), .in1(R4116));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4294 (.out1(R4295), .clock(clock), .in1(R4294));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4468 (.out1(R4469), .clock(clock), .in1(R4468));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4687 (.out1(R4688), .clock(clock), .in1(R4687));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4851 (.out1(R4852), .clock(clock), .in1(R4851));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5011 (.out1(R5012), .clock(clock), .in1(R5011));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5216 (.out1(R5217), .clock(clock), .in1(R5216));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5366 (.out1(R5367), .clock(clock), .in1(R5366));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5512 (.out1(R5513), .clock(clock), .in1(R5512));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5703 (.out1(R5704), .clock(clock), .in1(R5703));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5839 (.out1(R5840), .clock(clock), .in1(R5839));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5971 (.out1(R5972), .clock(clock), .in1(R5971));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6147 (.out1(R6148), .clock(clock), .in1(R6147));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6268 (.out1(R6269), .clock(clock), .in1(R6268));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6385 (.out1(R6386), .clock(clock), .in1(R6385));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6548 (.out1(R6549), .clock(clock), .in1(R6548));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6655 (.out1(R6656), .clock(clock), .in1(R6655));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6758 (.out1(R6759), .clock(clock), .in1(R6758));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6906 (.out1(R6907), .clock(clock), .in1(R6906));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6999 (.out1(R7000), .clock(clock), .in1(R6999));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7088 (.out1(R7089), .clock(clock), .in1(R7088));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7222 (.out1(R7223), .clock(clock), .in1(R7222));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7301 (.out1(R7302), .clock(clock), .in1(R7301));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7376 (.out1(R7377), .clock(clock), .in1(R7376));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7496 (.out1(R7497), .clock(clock), .in1(R7496));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7561 (.out1(R7562), .clock(clock), .in1(R7561));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7622 (.out1(R7623), .clock(clock), .in1(R7622));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7728 (.out1(R7729), .clock(clock), .in1(R7728));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7779 (.out1(R7780), .clock(clock), .in1(R7779));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7826 (.out1(R7827), .clock(clock), .in1(R7826));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7918 (.out1(R7919), .clock(clock), .in1(R7918));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7955 (.out1(R7956), .clock(clock), .in1(R7955));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7988 (.out1(R7989), .clock(clock), .in1(R7988));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8057 (.out1(R8058), .clock(clock), .in1(_1063));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8058 (.out1(R8059), .clock(clock), .in1(_1133));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8059 (.out1(R8060), .clock(clock), .in1(_1097));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8060 (.out1(R8061), .clock(clock), .in1(_1080));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1161 (.out1(_1098), .in1(R8060), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1144 (.out1(_1081), .in1(R8061), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op1197 (.out1(_1134), .in1(R8059), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1162 (.out1(_1099), .in1(_1081), .in2(_1098));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1127 (.out1(_1064), .in1(c112_popcnt_2654_D), .in2(R8058));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1198 (.out1(_1135), .in1(_1099), .in2(_1134));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op1199 (.out1(_1136), .in1(_1135), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2849 (.out1(R2850), .clock(clock), .in1(R2849));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3055 (.out1(R3056), .clock(clock), .in1(R3055));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3257 (.out1(R3258), .clock(clock), .in1(R3257));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3504 (.out1(R3505), .clock(clock), .in1(R3504));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3696 (.out1(R3697), .clock(clock), .in1(R3696));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3884 (.out1(R3885), .clock(clock), .in1(R3884));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4117 (.out1(R4118), .clock(clock), .in1(R4117));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4295 (.out1(R4296), .clock(clock), .in1(R4295));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4469 (.out1(R4470), .clock(clock), .in1(R4469));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4688 (.out1(R4689), .clock(clock), .in1(R4688));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4852 (.out1(R4853), .clock(clock), .in1(R4852));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5012 (.out1(R5013), .clock(clock), .in1(R5012));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5217 (.out1(R5218), .clock(clock), .in1(R5217));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5367 (.out1(R5368), .clock(clock), .in1(R5367));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5513 (.out1(R5514), .clock(clock), .in1(R5513));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5704 (.out1(R5705), .clock(clock), .in1(R5704));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5840 (.out1(R5841), .clock(clock), .in1(R5840));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5972 (.out1(R5973), .clock(clock), .in1(R5972));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6148 (.out1(R6149), .clock(clock), .in1(R6148));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6269 (.out1(R6270), .clock(clock), .in1(R6269));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6386 (.out1(R6387), .clock(clock), .in1(R6386));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6549 (.out1(R6550), .clock(clock), .in1(R6549));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6656 (.out1(R6657), .clock(clock), .in1(R6656));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6759 (.out1(R6760), .clock(clock), .in1(R6759));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6907 (.out1(R6908), .clock(clock), .in1(R6907));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7000 (.out1(R7001), .clock(clock), .in1(R7000));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7089 (.out1(R7090), .clock(clock), .in1(R7089));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7223 (.out1(R7224), .clock(clock), .in1(R7223));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7302 (.out1(R7303), .clock(clock), .in1(R7302));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7377 (.out1(R7378), .clock(clock), .in1(R7377));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7497 (.out1(R7498), .clock(clock), .in1(R7497));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7562 (.out1(R7563), .clock(clock), .in1(R7562));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7623 (.out1(R7624), .clock(clock), .in1(R7623));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7729 (.out1(R7730), .clock(clock), .in1(R7729));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7780 (.out1(R7781), .clock(clock), .in1(R7780));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7827 (.out1(R7828), .clock(clock), .in1(R7827));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7919 (.out1(R7920), .clock(clock), .in1(R7919));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7956 (.out1(R7957), .clock(clock), .in1(R7956));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7989 (.out1(R7990), .clock(clock), .in1(R7989));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8061 (.out1(R8062), .clock(clock), .in1(_1064));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8062 (.out1(R8063), .clock(clock), .in1(_1136));
  SRAM op1128 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1065),.ADR(R8062));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op1200 (.out1(_1137), .in1(R8063), .in2(57 'd 72340172838076673));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2850 (.out1(R2851), .clock(clock), .in1(R2850));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3056 (.out1(R3057), .clock(clock), .in1(R3056));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3258 (.out1(R3259), .clock(clock), .in1(R3258));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3505 (.out1(R3506), .clock(clock), .in1(R3505));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3697 (.out1(R3698), .clock(clock), .in1(R3697));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3885 (.out1(R3886), .clock(clock), .in1(R3885));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4118 (.out1(R4119), .clock(clock), .in1(R4118));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4296 (.out1(R4297), .clock(clock), .in1(R4296));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4470 (.out1(R4471), .clock(clock), .in1(R4470));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4689 (.out1(R4690), .clock(clock), .in1(R4689));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4853 (.out1(R4854), .clock(clock), .in1(R4853));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5013 (.out1(R5014), .clock(clock), .in1(R5013));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5218 (.out1(R5219), .clock(clock), .in1(R5218));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5368 (.out1(R5369), .clock(clock), .in1(R5368));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5514 (.out1(R5515), .clock(clock), .in1(R5514));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5705 (.out1(R5706), .clock(clock), .in1(R5705));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5841 (.out1(R5842), .clock(clock), .in1(R5841));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5973 (.out1(R5974), .clock(clock), .in1(R5973));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6149 (.out1(R6150), .clock(clock), .in1(R6149));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6270 (.out1(R6271), .clock(clock), .in1(R6270));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6387 (.out1(R6388), .clock(clock), .in1(R6387));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6550 (.out1(R6551), .clock(clock), .in1(R6550));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6657 (.out1(R6658), .clock(clock), .in1(R6657));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6760 (.out1(R6761), .clock(clock), .in1(R6760));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6908 (.out1(R6909), .clock(clock), .in1(R6908));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7001 (.out1(R7002), .clock(clock), .in1(R7001));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7090 (.out1(R7091), .clock(clock), .in1(R7090));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7224 (.out1(R7225), .clock(clock), .in1(R7224));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7303 (.out1(R7304), .clock(clock), .in1(R7303));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7378 (.out1(R7379), .clock(clock), .in1(R7378));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7498 (.out1(R7499), .clock(clock), .in1(R7498));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7563 (.out1(R7564), .clock(clock), .in1(R7563));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7624 (.out1(R7625), .clock(clock), .in1(R7624));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7730 (.out1(R7731), .clock(clock), .in1(R7730));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7781 (.out1(R7782), .clock(clock), .in1(R7781));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7828 (.out1(R7829), .clock(clock), .in1(R7828));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7920 (.out1(R7921), .clock(clock), .in1(R7920));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7957 (.out1(R7958), .clock(clock), .in1(R7957));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7990 (.out1(R7991), .clock(clock), .in1(R7990));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8063 (.out1(R8064), .clock(clock), .in1(_1065));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8064 (.out1(R8065), .clock(clock), .in1(_1137));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op1201 (.out1(_1138), .in1(R8065), .in2(6 'd 56));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1202 (.out1(_1139), .in1(_1138));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1203 (.out1(ck_idx_2655), .in1(R8064), .in2(_1139));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2851 (.out1(R2852), .clock(clock), .in1(R2851));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3057 (.out1(R3058), .clock(clock), .in1(R3057));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3259 (.out1(R3260), .clock(clock), .in1(R3259));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3506 (.out1(R3507), .clock(clock), .in1(R3506));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3698 (.out1(R3699), .clock(clock), .in1(R3698));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3886 (.out1(R3887), .clock(clock), .in1(R3886));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4119 (.out1(R4120), .clock(clock), .in1(R4119));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4297 (.out1(R4298), .clock(clock), .in1(R4297));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4471 (.out1(R4472), .clock(clock), .in1(R4471));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4690 (.out1(R4691), .clock(clock), .in1(R4690));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4854 (.out1(R4855), .clock(clock), .in1(R4854));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5014 (.out1(R5015), .clock(clock), .in1(R5014));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5219 (.out1(R5220), .clock(clock), .in1(R5219));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5369 (.out1(R5370), .clock(clock), .in1(R5369));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5515 (.out1(R5516), .clock(clock), .in1(R5515));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5706 (.out1(R5707), .clock(clock), .in1(R5706));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5842 (.out1(R5843), .clock(clock), .in1(R5842));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5974 (.out1(R5975), .clock(clock), .in1(R5974));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6150 (.out1(R6151), .clock(clock), .in1(R6150));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6271 (.out1(R6272), .clock(clock), .in1(R6271));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6388 (.out1(R6389), .clock(clock), .in1(R6388));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6551 (.out1(R6552), .clock(clock), .in1(R6551));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6658 (.out1(R6659), .clock(clock), .in1(R6658));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6761 (.out1(R6762), .clock(clock), .in1(R6761));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6909 (.out1(R6910), .clock(clock), .in1(R6909));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7002 (.out1(R7003), .clock(clock), .in1(R7002));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7091 (.out1(R7092), .clock(clock), .in1(R7091));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7225 (.out1(R7226), .clock(clock), .in1(R7225));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7304 (.out1(R7305), .clock(clock), .in1(R7304));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7379 (.out1(R7380), .clock(clock), .in1(R7379));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7499 (.out1(R7500), .clock(clock), .in1(R7499));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7564 (.out1(R7565), .clock(clock), .in1(R7564));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7625 (.out1(R7626), .clock(clock), .in1(R7625));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7731 (.out1(R7732), .clock(clock), .in1(R7731));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7782 (.out1(R7783), .clock(clock), .in1(R7782));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7829 (.out1(R7830), .clock(clock), .in1(R7829));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7921 (.out1(R7922), .clock(clock), .in1(R7921));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7958 (.out1(R7959), .clock(clock), .in1(R7958));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7991 (.out1(R7992), .clock(clock), .in1(R7991));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8065 (.out1(R8066), .clock(clock), .in1(ck_idx_2655));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(4), .BITSIZE_out1(32), .PRECISION(32)) op1204 (.out1(_1140), .in1(R8066), .in2(4 'd 8));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(4), .BITSIZE_out1(64), .PRECISION(64)) op1205 (.out1(_1141), .in1(ip2_2595_D), .in2(4 'd 8));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2852 (.out1(R2853), .clock(clock), .in1(R2852));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3058 (.out1(R3059), .clock(clock), .in1(R3058));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3260 (.out1(R3261), .clock(clock), .in1(R3260));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3507 (.out1(R3508), .clock(clock), .in1(R3507));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3699 (.out1(R3700), .clock(clock), .in1(R3699));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3887 (.out1(R3888), .clock(clock), .in1(R3887));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4120 (.out1(R4121), .clock(clock), .in1(R4120));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4298 (.out1(R4299), .clock(clock), .in1(R4298));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4472 (.out1(R4473), .clock(clock), .in1(R4472));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4691 (.out1(R4692), .clock(clock), .in1(R4691));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4855 (.out1(R4856), .clock(clock), .in1(R4855));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5015 (.out1(R5016), .clock(clock), .in1(R5015));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5220 (.out1(R5221), .clock(clock), .in1(R5220));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5370 (.out1(R5371), .clock(clock), .in1(R5370));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5516 (.out1(R5517), .clock(clock), .in1(R5516));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5707 (.out1(R5708), .clock(clock), .in1(R5707));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5843 (.out1(R5844), .clock(clock), .in1(R5843));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5975 (.out1(R5976), .clock(clock), .in1(R5975));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6151 (.out1(R6152), .clock(clock), .in1(R6151));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6272 (.out1(R6273), .clock(clock), .in1(R6272));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6389 (.out1(R6390), .clock(clock), .in1(R6389));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6552 (.out1(R6553), .clock(clock), .in1(R6552));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6659 (.out1(R6660), .clock(clock), .in1(R6659));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6762 (.out1(R6763), .clock(clock), .in1(R6762));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6910 (.out1(R6911), .clock(clock), .in1(R6910));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7003 (.out1(R7004), .clock(clock), .in1(R7003));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7092 (.out1(R7093), .clock(clock), .in1(R7092));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7226 (.out1(R7227), .clock(clock), .in1(R7226));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7305 (.out1(R7306), .clock(clock), .in1(R7305));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7380 (.out1(R7381), .clock(clock), .in1(R7380));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7500 (.out1(R7501), .clock(clock), .in1(R7500));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7565 (.out1(R7566), .clock(clock), .in1(R7565));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7626 (.out1(R7627), .clock(clock), .in1(R7626));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7732 (.out1(R7733), .clock(clock), .in1(R7732));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7783 (.out1(R7784), .clock(clock), .in1(R7783));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7830 (.out1(R7831), .clock(clock), .in1(R7830));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7922 (.out1(R7923), .clock(clock), .in1(R7922));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7959 (.out1(R7960), .clock(clock), .in1(R7959));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7992 (.out1(R7993), .clock(clock), .in1(R7992));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8066 (.out1(R8067), .clock(clock), .in1(_1140));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8067 (.out1(R8068), .clock(clock), .in1(_1141));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1206 (.out1(_1142), .in1(R8068));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(8), .BITSIZE_out1(32)) op1207 (.out1(_1143), .in1(_1142), .in2(8 'd 255));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1208 (.out1(idx_sail_2656), .in1(R8067), .in2(_1143));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(3), .BITSIZE_out1(32), .PRECISION(32)) op1209 (.out1(idx_2657), .in1(idx_sail_2656), .in2(3 'd 6));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2853 (.out1(R2854), .clock(clock), .in1(R2853));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3059 (.out1(R3060), .clock(clock), .in1(R3059));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3261 (.out1(R3262), .clock(clock), .in1(R3261));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3508 (.out1(R3509), .clock(clock), .in1(R3508));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3700 (.out1(R3701), .clock(clock), .in1(R3700));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3888 (.out1(R3889), .clock(clock), .in1(R3888));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4121 (.out1(R4122), .clock(clock), .in1(R4121));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4299 (.out1(R4300), .clock(clock), .in1(R4299));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4473 (.out1(R4474), .clock(clock), .in1(R4473));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4692 (.out1(R4693), .clock(clock), .in1(R4692));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4856 (.out1(R4857), .clock(clock), .in1(R4856));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5016 (.out1(R5017), .clock(clock), .in1(R5016));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5221 (.out1(R5222), .clock(clock), .in1(R5221));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5371 (.out1(R5372), .clock(clock), .in1(R5371));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5517 (.out1(R5518), .clock(clock), .in1(R5517));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5708 (.out1(R5709), .clock(clock), .in1(R5708));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5844 (.out1(R5845), .clock(clock), .in1(R5844));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5976 (.out1(R5977), .clock(clock), .in1(R5976));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6152 (.out1(R6153), .clock(clock), .in1(R6152));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6273 (.out1(R6274), .clock(clock), .in1(R6273));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6390 (.out1(R6391), .clock(clock), .in1(R6390));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6553 (.out1(R6554), .clock(clock), .in1(R6553));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6660 (.out1(R6661), .clock(clock), .in1(R6660));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6763 (.out1(R6764), .clock(clock), .in1(R6763));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6911 (.out1(R6912), .clock(clock), .in1(R6911));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7004 (.out1(R7005), .clock(clock), .in1(R7004));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7093 (.out1(R7094), .clock(clock), .in1(R7093));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7227 (.out1(R7228), .clock(clock), .in1(R7227));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7306 (.out1(R7307), .clock(clock), .in1(R7306));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7381 (.out1(R7382), .clock(clock), .in1(R7381));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7501 (.out1(R7502), .clock(clock), .in1(R7501));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7566 (.out1(R7567), .clock(clock), .in1(R7566));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7627 (.out1(R7628), .clock(clock), .in1(R7627));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7733 (.out1(R7734), .clock(clock), .in1(R7733));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7784 (.out1(R7785), .clock(clock), .in1(R7784));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7831 (.out1(R7832), .clock(clock), .in1(R7831));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7923 (.out1(R7924), .clock(clock), .in1(R7923));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7960 (.out1(R7961), .clock(clock), .in1(R7960));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7993 (.out1(R7994), .clock(clock), .in1(R7993));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8068 (.out1(R8069), .clock(clock), .in1(idx_sail_2656));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8071 (.out1(R8072), .clock(clock), .in1(idx_2657));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1211 (.out1(_1144), .in1(R8072));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1212 (.out1(_1145), .in1(_1144), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2854 (.out1(R2855), .clock(clock), .in1(R2854));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3060 (.out1(R3061), .clock(clock), .in1(R3060));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3262 (.out1(R3263), .clock(clock), .in1(R3262));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3509 (.out1(R3510), .clock(clock), .in1(R3509));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3701 (.out1(R3702), .clock(clock), .in1(R3701));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3889 (.out1(R3890), .clock(clock), .in1(R3889));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4122 (.out1(R4123), .clock(clock), .in1(R4122));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4300 (.out1(R4301), .clock(clock), .in1(R4300));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4474 (.out1(R4475), .clock(clock), .in1(R4474));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4693 (.out1(R4694), .clock(clock), .in1(R4693));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4857 (.out1(R4858), .clock(clock), .in1(R4857));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5017 (.out1(R5018), .clock(clock), .in1(R5017));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5222 (.out1(R5223), .clock(clock), .in1(R5222));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5372 (.out1(R5373), .clock(clock), .in1(R5372));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5518 (.out1(R5519), .clock(clock), .in1(R5518));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5709 (.out1(R5710), .clock(clock), .in1(R5709));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5845 (.out1(R5846), .clock(clock), .in1(R5845));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5977 (.out1(R5978), .clock(clock), .in1(R5977));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6153 (.out1(R6154), .clock(clock), .in1(R6153));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6274 (.out1(R6275), .clock(clock), .in1(R6274));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6391 (.out1(R6392), .clock(clock), .in1(R6391));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6554 (.out1(R6555), .clock(clock), .in1(R6554));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6661 (.out1(R6662), .clock(clock), .in1(R6661));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6764 (.out1(R6765), .clock(clock), .in1(R6764));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6912 (.out1(R6913), .clock(clock), .in1(R6912));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7005 (.out1(R7006), .clock(clock), .in1(R7005));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7094 (.out1(R7095), .clock(clock), .in1(R7094));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7228 (.out1(R7229), .clock(clock), .in1(R7228));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7307 (.out1(R7308), .clock(clock), .in1(R7307));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7382 (.out1(R7383), .clock(clock), .in1(R7382));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7502 (.out1(R7503), .clock(clock), .in1(R7502));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7567 (.out1(R7568), .clock(clock), .in1(R7567));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7628 (.out1(R7629), .clock(clock), .in1(R7628));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7734 (.out1(R7735), .clock(clock), .in1(R7734));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7785 (.out1(R7786), .clock(clock), .in1(R7785));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7832 (.out1(R7833), .clock(clock), .in1(R7832));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7924 (.out1(R7925), .clock(clock), .in1(R7924));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7961 (.out1(R7962), .clock(clock), .in1(R7961));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7994 (.out1(R7995), .clock(clock), .in1(R7994));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8069 (.out1(R8070), .clock(clock), .in1(R8069));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8072 (.out1(R8073), .clock(clock), .in1(R8072));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8094 (.out1(R8095), .clock(clock), .in1(_1145));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1213 (.out1(_1146), .in1(c120_bitmap_2659_D), .in2(R8095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2855 (.out1(R2856), .clock(clock), .in1(R2855));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3061 (.out1(R3062), .clock(clock), .in1(R3061));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3263 (.out1(R3264), .clock(clock), .in1(R3263));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3510 (.out1(R3511), .clock(clock), .in1(R3510));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3702 (.out1(R3703), .clock(clock), .in1(R3702));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3890 (.out1(R3891), .clock(clock), .in1(R3890));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4123 (.out1(R4124), .clock(clock), .in1(R4123));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4301 (.out1(R4302), .clock(clock), .in1(R4301));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4475 (.out1(R4476), .clock(clock), .in1(R4475));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4694 (.out1(R4695), .clock(clock), .in1(R4694));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4858 (.out1(R4859), .clock(clock), .in1(R4858));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5018 (.out1(R5019), .clock(clock), .in1(R5018));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5223 (.out1(R5224), .clock(clock), .in1(R5223));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5373 (.out1(R5374), .clock(clock), .in1(R5373));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5519 (.out1(R5520), .clock(clock), .in1(R5519));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5710 (.out1(R5711), .clock(clock), .in1(R5710));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5846 (.out1(R5847), .clock(clock), .in1(R5846));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5978 (.out1(R5979), .clock(clock), .in1(R5978));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6154 (.out1(R6155), .clock(clock), .in1(R6154));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6275 (.out1(R6276), .clock(clock), .in1(R6275));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6392 (.out1(R6393), .clock(clock), .in1(R6392));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6555 (.out1(R6556), .clock(clock), .in1(R6555));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6662 (.out1(R6663), .clock(clock), .in1(R6662));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6765 (.out1(R6766), .clock(clock), .in1(R6765));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6913 (.out1(R6914), .clock(clock), .in1(R6913));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7006 (.out1(R7007), .clock(clock), .in1(R7006));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7095 (.out1(R7096), .clock(clock), .in1(R7095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7229 (.out1(R7230), .clock(clock), .in1(R7229));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7308 (.out1(R7309), .clock(clock), .in1(R7308));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7383 (.out1(R7384), .clock(clock), .in1(R7383));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7503 (.out1(R7504), .clock(clock), .in1(R7503));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7568 (.out1(R7569), .clock(clock), .in1(R7568));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7629 (.out1(R7630), .clock(clock), .in1(R7629));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7735 (.out1(R7736), .clock(clock), .in1(R7735));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7786 (.out1(R7787), .clock(clock), .in1(R7786));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7833 (.out1(R7834), .clock(clock), .in1(R7833));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7925 (.out1(R7926), .clock(clock), .in1(R7925));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7962 (.out1(R7963), .clock(clock), .in1(R7962));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7995 (.out1(R7996), .clock(clock), .in1(R7995));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8070 (.out1(R8071), .clock(clock), .in1(R8070));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8073 (.out1(R8074), .clock(clock), .in1(R8073));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8095 (.out1(R8096), .clock(clock), .in1(_1146));
  SRAM op1214 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1147),.ADR(R8096));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op1210 (.out1(off_2658), .in1(R8071), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1215 (.out1(_1148), .in1(64 'd 9223372036854775808), .in2(off_2658));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2856 (.out1(R2857), .clock(clock), .in1(R2856));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3062 (.out1(R3063), .clock(clock), .in1(R3062));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3264 (.out1(R3265), .clock(clock), .in1(R3264));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3511 (.out1(R3512), .clock(clock), .in1(R3511));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3703 (.out1(R3704), .clock(clock), .in1(R3703));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3891 (.out1(R3892), .clock(clock), .in1(R3891));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4124 (.out1(R4125), .clock(clock), .in1(R4124));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4302 (.out1(R4303), .clock(clock), .in1(R4302));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4476 (.out1(R4477), .clock(clock), .in1(R4476));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4695 (.out1(R4696), .clock(clock), .in1(R4695));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4859 (.out1(R4860), .clock(clock), .in1(R4859));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5019 (.out1(R5020), .clock(clock), .in1(R5019));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5224 (.out1(R5225), .clock(clock), .in1(R5224));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5374 (.out1(R5375), .clock(clock), .in1(R5374));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5520 (.out1(R5521), .clock(clock), .in1(R5520));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5711 (.out1(R5712), .clock(clock), .in1(R5711));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5847 (.out1(R5848), .clock(clock), .in1(R5847));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5979 (.out1(R5980), .clock(clock), .in1(R5979));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6155 (.out1(R6156), .clock(clock), .in1(R6155));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6276 (.out1(R6277), .clock(clock), .in1(R6276));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6393 (.out1(R6394), .clock(clock), .in1(R6393));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6556 (.out1(R6557), .clock(clock), .in1(R6556));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6663 (.out1(R6664), .clock(clock), .in1(R6663));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6766 (.out1(R6767), .clock(clock), .in1(R6766));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6914 (.out1(R6915), .clock(clock), .in1(R6914));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7007 (.out1(R7008), .clock(clock), .in1(R7007));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7096 (.out1(R7097), .clock(clock), .in1(R7096));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7230 (.out1(R7231), .clock(clock), .in1(R7230));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7309 (.out1(R7310), .clock(clock), .in1(R7309));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7384 (.out1(R7385), .clock(clock), .in1(R7384));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7504 (.out1(R7505), .clock(clock), .in1(R7504));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7569 (.out1(R7570), .clock(clock), .in1(R7569));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7630 (.out1(R7631), .clock(clock), .in1(R7630));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7736 (.out1(R7737), .clock(clock), .in1(R7736));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7787 (.out1(R7788), .clock(clock), .in1(R7787));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7834 (.out1(R7835), .clock(clock), .in1(R7834));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7926 (.out1(R7927), .clock(clock), .in1(R7926));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7963 (.out1(R7964), .clock(clock), .in1(R7963));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7996 (.out1(R7997), .clock(clock), .in1(R7996));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8074 (.out1(R8075), .clock(clock), .in1(R8074));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8096 (.out1(R8097), .clock(clock), .in1(_1147));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8097 (.out1(R8098), .clock(clock), .in1(off_2658));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8116 (.out1(R8117), .clock(clock), .in1(_1148));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1216 (.out1(_1149), .in1(R8097), .in2(R8117));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op1217 (.out1(ifout1217), .in1(_1149), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1278 (.out1(_1210), .in1(R8075));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1279 (.out1(_1211), .in1(_1210), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2857 (.out1(R2858), .clock(clock), .in1(R2857));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3063 (.out1(R3064), .clock(clock), .in1(R3063));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3265 (.out1(R3266), .clock(clock), .in1(R3265));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3512 (.out1(R3513), .clock(clock), .in1(R3512));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3704 (.out1(R3705), .clock(clock), .in1(R3704));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3892 (.out1(R3893), .clock(clock), .in1(R3892));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4125 (.out1(R4126), .clock(clock), .in1(R4125));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4303 (.out1(R4304), .clock(clock), .in1(R4303));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4477 (.out1(R4478), .clock(clock), .in1(R4477));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4696 (.out1(R4697), .clock(clock), .in1(R4696));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4860 (.out1(R4861), .clock(clock), .in1(R4860));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5020 (.out1(R5021), .clock(clock), .in1(R5020));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5225 (.out1(R5226), .clock(clock), .in1(R5225));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5375 (.out1(R5376), .clock(clock), .in1(R5375));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5521 (.out1(R5522), .clock(clock), .in1(R5521));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5712 (.out1(R5713), .clock(clock), .in1(R5712));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5848 (.out1(R5849), .clock(clock), .in1(R5848));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5980 (.out1(R5981), .clock(clock), .in1(R5980));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6156 (.out1(R6157), .clock(clock), .in1(R6156));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6277 (.out1(R6278), .clock(clock), .in1(R6277));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6394 (.out1(R6395), .clock(clock), .in1(R6394));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6557 (.out1(R6558), .clock(clock), .in1(R6557));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6664 (.out1(R6665), .clock(clock), .in1(R6664));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6767 (.out1(R6768), .clock(clock), .in1(R6767));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6915 (.out1(R6916), .clock(clock), .in1(R6915));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7008 (.out1(R7009), .clock(clock), .in1(R7008));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7097 (.out1(R7098), .clock(clock), .in1(R7097));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7231 (.out1(R7232), .clock(clock), .in1(R7231));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7310 (.out1(R7311), .clock(clock), .in1(R7310));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7385 (.out1(R7386), .clock(clock), .in1(R7385));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7505 (.out1(R7506), .clock(clock), .in1(R7505));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7570 (.out1(R7571), .clock(clock), .in1(R7570));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7631 (.out1(R7632), .clock(clock), .in1(R7631));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7737 (.out1(R7738), .clock(clock), .in1(R7737));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7788 (.out1(R7789), .clock(clock), .in1(R7788));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7835 (.out1(R7836), .clock(clock), .in1(R7835));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7927 (.out1(R7928), .clock(clock), .in1(R7927));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7964 (.out1(R7965), .clock(clock), .in1(R7964));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7997 (.out1(R7998), .clock(clock), .in1(R7997));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8075 (.out1(R8076), .clock(clock), .in1(R8075));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8098 (.out1(R8099), .clock(clock), .in1(R8098));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8117 (.out1(R8118), .clock(clock), .in1(ifout1217));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8142 (.out1(R8143), .clock(clock), .in1(_1211));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1272 (.out1(_1204), .in1(R8076));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1262 (.out1(_1194), .in1(R8076));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1256 (.out1(_1188), .in1(R8076));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1244 (.out1(_1176), .in1(R8076));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1238 (.out1(_1170), .in1(R8076));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1228 (.out1(_1160), .in1(R8076));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1273 (.out1(_1205), .in1(_1204), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1263 (.out1(_1195), .in1(_1194), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1257 (.out1(_1189), .in1(_1188), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1245 (.out1(_1177), .in1(_1176), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1239 (.out1(_1171), .in1(_1170), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1229 (.out1(_1161), .in1(_1160), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1280 (.out1(_1212), .in1(c120_bitmap_2659_D), .in2(R8143));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2858 (.out1(R2859), .clock(clock), .in1(R2858));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3064 (.out1(R3065), .clock(clock), .in1(R3064));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3266 (.out1(R3267), .clock(clock), .in1(R3266));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3513 (.out1(R3514), .clock(clock), .in1(R3513));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3705 (.out1(R3706), .clock(clock), .in1(R3705));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3893 (.out1(R3894), .clock(clock), .in1(R3893));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4126 (.out1(R4127), .clock(clock), .in1(R4126));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4304 (.out1(R4305), .clock(clock), .in1(R4304));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4478 (.out1(R4479), .clock(clock), .in1(R4478));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4697 (.out1(R4698), .clock(clock), .in1(R4697));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4861 (.out1(R4862), .clock(clock), .in1(R4861));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5021 (.out1(R5022), .clock(clock), .in1(R5021));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5226 (.out1(R5227), .clock(clock), .in1(R5226));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5376 (.out1(R5377), .clock(clock), .in1(R5376));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5522 (.out1(R5523), .clock(clock), .in1(R5522));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5713 (.out1(R5714), .clock(clock), .in1(R5713));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5849 (.out1(R5850), .clock(clock), .in1(R5849));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5981 (.out1(R5982), .clock(clock), .in1(R5981));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6157 (.out1(R6158), .clock(clock), .in1(R6157));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6278 (.out1(R6279), .clock(clock), .in1(R6278));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6395 (.out1(R6396), .clock(clock), .in1(R6395));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6558 (.out1(R6559), .clock(clock), .in1(R6558));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6665 (.out1(R6666), .clock(clock), .in1(R6665));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6768 (.out1(R6769), .clock(clock), .in1(R6768));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6916 (.out1(R6917), .clock(clock), .in1(R6916));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7009 (.out1(R7010), .clock(clock), .in1(R7009));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7098 (.out1(R7099), .clock(clock), .in1(R7098));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7232 (.out1(R7233), .clock(clock), .in1(R7232));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7311 (.out1(R7312), .clock(clock), .in1(R7311));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7386 (.out1(R7387), .clock(clock), .in1(R7386));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7506 (.out1(R7507), .clock(clock), .in1(R7506));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7571 (.out1(R7572), .clock(clock), .in1(R7571));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7632 (.out1(R7633), .clock(clock), .in1(R7632));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7738 (.out1(R7739), .clock(clock), .in1(R7738));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7789 (.out1(R7790), .clock(clock), .in1(R7789));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7836 (.out1(R7837), .clock(clock), .in1(R7836));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7928 (.out1(R7929), .clock(clock), .in1(R7928));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7965 (.out1(R7966), .clock(clock), .in1(R7965));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7998 (.out1(R7999), .clock(clock), .in1(R7998));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8076 (.out1(R8077), .clock(clock), .in1(R8076));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8099 (.out1(R8100), .clock(clock), .in1(R8099));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8118 (.out1(R8119), .clock(clock), .in1(R8118));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8143 (.out1(R8144), .clock(clock), .in1(_1205));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8144 (.out1(R8145), .clock(clock), .in1(_1195));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8145 (.out1(R8146), .clock(clock), .in1(_1189));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8146 (.out1(R8147), .clock(clock), .in1(_1177));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8147 (.out1(R8148), .clock(clock), .in1(_1171));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8148 (.out1(R8149), .clock(clock), .in1(_1161));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8149 (.out1(R8150), .clock(clock), .in1(_1212));
  SRAM op1281 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1213),.ADR(R8150));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1222 (.out1(_1154), .in1(R8077));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1223 (.out1(_1155), .in1(_1154), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1274 (.out1(_1206), .in1(c120_bitmap_2659_D), .in2(R8144));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1264 (.out1(_1196), .in1(c120_bitmap_2659_D), .in2(R8145));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1258 (.out1(_1190), .in1(c120_bitmap_2659_D), .in2(R8146));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1246 (.out1(_1178), .in1(c120_bitmap_2659_D), .in2(R8147));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1240 (.out1(_1172), .in1(c120_bitmap_2659_D), .in2(R8148));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1230 (.out1(_1162), .in1(c120_bitmap_2659_D), .in2(R8149));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2859 (.out1(R2860), .clock(clock), .in1(R2859));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3065 (.out1(R3066), .clock(clock), .in1(R3065));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3267 (.out1(R3268), .clock(clock), .in1(R3267));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3514 (.out1(R3515), .clock(clock), .in1(R3514));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3706 (.out1(R3707), .clock(clock), .in1(R3706));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3894 (.out1(R3895), .clock(clock), .in1(R3894));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4127 (.out1(R4128), .clock(clock), .in1(R4127));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4305 (.out1(R4306), .clock(clock), .in1(R4305));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4479 (.out1(R4480), .clock(clock), .in1(R4479));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4698 (.out1(R4699), .clock(clock), .in1(R4698));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4862 (.out1(R4863), .clock(clock), .in1(R4862));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5022 (.out1(R5023), .clock(clock), .in1(R5022));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5227 (.out1(R5228), .clock(clock), .in1(R5227));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5377 (.out1(R5378), .clock(clock), .in1(R5377));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5523 (.out1(R5524), .clock(clock), .in1(R5523));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5714 (.out1(R5715), .clock(clock), .in1(R5714));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5850 (.out1(R5851), .clock(clock), .in1(R5850));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5982 (.out1(R5983), .clock(clock), .in1(R5982));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6158 (.out1(R6159), .clock(clock), .in1(R6158));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6279 (.out1(R6280), .clock(clock), .in1(R6279));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6396 (.out1(R6397), .clock(clock), .in1(R6396));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6559 (.out1(R6560), .clock(clock), .in1(R6559));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6666 (.out1(R6667), .clock(clock), .in1(R6666));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6769 (.out1(R6770), .clock(clock), .in1(R6769));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6917 (.out1(R6918), .clock(clock), .in1(R6917));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7010 (.out1(R7011), .clock(clock), .in1(R7010));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7099 (.out1(R7100), .clock(clock), .in1(R7099));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7233 (.out1(R7234), .clock(clock), .in1(R7233));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7312 (.out1(R7313), .clock(clock), .in1(R7312));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7387 (.out1(R7388), .clock(clock), .in1(R7387));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7507 (.out1(R7508), .clock(clock), .in1(R7507));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7572 (.out1(R7573), .clock(clock), .in1(R7572));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7633 (.out1(R7634), .clock(clock), .in1(R7633));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7739 (.out1(R7740), .clock(clock), .in1(R7739));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7790 (.out1(R7791), .clock(clock), .in1(R7790));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7837 (.out1(R7838), .clock(clock), .in1(R7837));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7929 (.out1(R7930), .clock(clock), .in1(R7929));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7966 (.out1(R7967), .clock(clock), .in1(R7966));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7999 (.out1(R8000), .clock(clock), .in1(R7999));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8077 (.out1(R8078), .clock(clock), .in1(R8077));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8100 (.out1(R8101), .clock(clock), .in1(R8100));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8119 (.out1(R8120), .clock(clock), .in1(R8119));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8150 (.out1(R8151), .clock(clock), .in1(_1213));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8151 (.out1(R8152), .clock(clock), .in1(_1155));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8152 (.out1(R8153), .clock(clock), .in1(_1206));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8153 (.out1(R8154), .clock(clock), .in1(_1196));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8154 (.out1(R8155), .clock(clock), .in1(_1190));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8155 (.out1(R8156), .clock(clock), .in1(_1178));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8156 (.out1(R8157), .clock(clock), .in1(_1172));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8157 (.out1(R8158), .clock(clock), .in1(_1162));
  SRAM op1275 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1207),.ADR(R8153));
  SRAM op1265 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1197),.ADR(R8154));
  SRAM op1259 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1191),.ADR(R8155));
  SRAM op1247 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1179),.ADR(R8156));
  SRAM op1241 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1173),.ADR(R8157));
  SRAM op1231 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1163),.ADR(R8158));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1282 (.out1(_1214), .in1(7 'd 64), .in2(R8101));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1224 (.out1(_1156), .in1(c120_bitmap_2659_D), .in2(R8152));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1283 (.out1(_1215), .in1(R8151), .in2(_1214));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1276 (.out1(_1208), .in1(7 'd 64), .in2(R8101));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1266 (.out1(_1198), .in1(7 'd 64), .in2(R8101));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1248 (.out1(_1180), .in1(7 'd 64), .in2(R8101));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2860 (.out1(R2861), .clock(clock), .in1(R2860));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3066 (.out1(R3067), .clock(clock), .in1(R3066));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3268 (.out1(R3269), .clock(clock), .in1(R3268));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3515 (.out1(R3516), .clock(clock), .in1(R3515));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3707 (.out1(R3708), .clock(clock), .in1(R3707));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3895 (.out1(R3896), .clock(clock), .in1(R3895));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4128 (.out1(R4129), .clock(clock), .in1(R4128));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4306 (.out1(R4307), .clock(clock), .in1(R4306));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4480 (.out1(R4481), .clock(clock), .in1(R4480));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4699 (.out1(R4700), .clock(clock), .in1(R4699));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4863 (.out1(R4864), .clock(clock), .in1(R4863));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5023 (.out1(R5024), .clock(clock), .in1(R5023));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5228 (.out1(R5229), .clock(clock), .in1(R5228));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5378 (.out1(R5379), .clock(clock), .in1(R5378));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5524 (.out1(R5525), .clock(clock), .in1(R5524));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5715 (.out1(R5716), .clock(clock), .in1(R5715));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5851 (.out1(R5852), .clock(clock), .in1(R5851));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5983 (.out1(R5984), .clock(clock), .in1(R5983));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6159 (.out1(R6160), .clock(clock), .in1(R6159));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6280 (.out1(R6281), .clock(clock), .in1(R6280));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6397 (.out1(R6398), .clock(clock), .in1(R6397));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6560 (.out1(R6561), .clock(clock), .in1(R6560));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6667 (.out1(R6668), .clock(clock), .in1(R6667));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6770 (.out1(R6771), .clock(clock), .in1(R6770));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6918 (.out1(R6919), .clock(clock), .in1(R6918));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7011 (.out1(R7012), .clock(clock), .in1(R7011));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7100 (.out1(R7101), .clock(clock), .in1(R7100));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7234 (.out1(R7235), .clock(clock), .in1(R7234));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7313 (.out1(R7314), .clock(clock), .in1(R7313));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7388 (.out1(R7389), .clock(clock), .in1(R7388));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7508 (.out1(R7509), .clock(clock), .in1(R7508));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7573 (.out1(R7574), .clock(clock), .in1(R7573));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7634 (.out1(R7635), .clock(clock), .in1(R7634));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7740 (.out1(R7741), .clock(clock), .in1(R7740));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7791 (.out1(R7792), .clock(clock), .in1(R7791));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7838 (.out1(R7839), .clock(clock), .in1(R7838));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7930 (.out1(R7931), .clock(clock), .in1(R7930));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7967 (.out1(R7968), .clock(clock), .in1(R7967));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8000 (.out1(R8001), .clock(clock), .in1(R8000));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8078 (.out1(R8079), .clock(clock), .in1(R8078));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8101 (.out1(R8102), .clock(clock), .in1(R8101));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8120 (.out1(R8121), .clock(clock), .in1(R8120));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8158 (.out1(R8159), .clock(clock), .in1(_1207));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8159 (.out1(R8160), .clock(clock), .in1(_1197));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8160 (.out1(R8161), .clock(clock), .in1(_1191));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8161 (.out1(R8162), .clock(clock), .in1(_1179));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8162 (.out1(R8163), .clock(clock), .in1(_1173));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8163 (.out1(R8164), .clock(clock), .in1(_1163));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8164 (.out1(R8165), .clock(clock), .in1(_1156));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8165 (.out1(R8166), .clock(clock), .in1(_1215));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8166 (.out1(R8167), .clock(clock), .in1(_1208));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8167 (.out1(R8168), .clock(clock), .in1(_1198));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8168 (.out1(R8169), .clock(clock), .in1(_1180));
  SRAM op1225 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1157),.ADR(R8165));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1284 (.out1(_1216), .in1(R8166), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1277 (.out1(_1209), .in1(R8159), .in2(R8167));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1267 (.out1(_1199), .in1(R8160), .in2(R8168));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1260 (.out1(_1192), .in1(7 'd 64), .in2(R8102));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1249 (.out1(_1181), .in1(R8162), .in2(R8169));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1242 (.out1(_1174), .in1(7 'd 64), .in2(R8102));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1232 (.out1(_1164), .in1(7 'd 64), .in2(R8102));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1285 (.out1(_1217), .in1(_1216), .in2(63 'd 6148914691236517205));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1286 (.out1(_1218), .in1(_1209), .in2(_1217));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1268 (.out1(_1200), .in1(_1199), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1261 (.out1(_1193), .in1(R8161), .in2(_1192));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1250 (.out1(_1182), .in1(_1181), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1243 (.out1(_1175), .in1(R8163), .in2(_1174));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1233 (.out1(_1165), .in1(R8164), .in2(_1164));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1226 (.out1(_1158), .in1(7 'd 64), .in2(R8102));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2861 (.out1(R2862), .clock(clock), .in1(R2861));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3067 (.out1(R3068), .clock(clock), .in1(R3067));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3269 (.out1(R3270), .clock(clock), .in1(R3269));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3516 (.out1(R3517), .clock(clock), .in1(R3516));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3708 (.out1(R3709), .clock(clock), .in1(R3708));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3896 (.out1(R3897), .clock(clock), .in1(R3896));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4129 (.out1(R4130), .clock(clock), .in1(R4129));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4307 (.out1(R4308), .clock(clock), .in1(R4307));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4481 (.out1(R4482), .clock(clock), .in1(R4481));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4700 (.out1(R4701), .clock(clock), .in1(R4700));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4864 (.out1(R4865), .clock(clock), .in1(R4864));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5024 (.out1(R5025), .clock(clock), .in1(R5024));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5229 (.out1(R5230), .clock(clock), .in1(R5229));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5379 (.out1(R5380), .clock(clock), .in1(R5379));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5525 (.out1(R5526), .clock(clock), .in1(R5525));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5716 (.out1(R5717), .clock(clock), .in1(R5716));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5852 (.out1(R5853), .clock(clock), .in1(R5852));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5984 (.out1(R5985), .clock(clock), .in1(R5984));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6160 (.out1(R6161), .clock(clock), .in1(R6160));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6281 (.out1(R6282), .clock(clock), .in1(R6281));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6398 (.out1(R6399), .clock(clock), .in1(R6398));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6561 (.out1(R6562), .clock(clock), .in1(R6561));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6668 (.out1(R6669), .clock(clock), .in1(R6668));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6771 (.out1(R6772), .clock(clock), .in1(R6771));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6919 (.out1(R6920), .clock(clock), .in1(R6919));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7012 (.out1(R7013), .clock(clock), .in1(R7012));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7101 (.out1(R7102), .clock(clock), .in1(R7101));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7235 (.out1(R7236), .clock(clock), .in1(R7235));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7314 (.out1(R7315), .clock(clock), .in1(R7314));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7389 (.out1(R7390), .clock(clock), .in1(R7389));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7509 (.out1(R7510), .clock(clock), .in1(R7509));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7574 (.out1(R7575), .clock(clock), .in1(R7574));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7635 (.out1(R7636), .clock(clock), .in1(R7635));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7741 (.out1(R7742), .clock(clock), .in1(R7741));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7792 (.out1(R7793), .clock(clock), .in1(R7792));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7839 (.out1(R7840), .clock(clock), .in1(R7839));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7931 (.out1(R7932), .clock(clock), .in1(R7931));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7968 (.out1(R7969), .clock(clock), .in1(R7968));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8001 (.out1(R8002), .clock(clock), .in1(R8001));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8079 (.out1(R8080), .clock(clock), .in1(R8079));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8102 (.out1(R8103), .clock(clock), .in1(R8102));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8121 (.out1(R8122), .clock(clock), .in1(R8121));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8169 (.out1(R8170), .clock(clock), .in1(_1157));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8170 (.out1(R8171), .clock(clock), .in1(_1218));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8171 (.out1(R8172), .clock(clock), .in1(_1200));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8172 (.out1(R8173), .clock(clock), .in1(_1193));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8173 (.out1(R8174), .clock(clock), .in1(_1182));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8174 (.out1(R8175), .clock(clock), .in1(_1175));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8175 (.out1(R8176), .clock(clock), .in1(_1165));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8176 (.out1(R8177), .clock(clock), .in1(_1158));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1218 (.out1(_1150), .in1(R8080));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1269 (.out1(_1201), .in1(R8172), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1287 (.out1(_1219), .in1(R8171), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1270 (.out1(_1202), .in1(R8173), .in2(_1201));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1251 (.out1(_1183), .in1(R8174), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1234 (.out1(_1166), .in1(R8176), .in2(1 'd 1));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1252 (.out1(_1184), .in1(R8175), .in2(_1183));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1227 (.out1(_1159), .in1(R8170), .in2(R8177));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1219 (.out1(_1151), .in1(_1150), .in2(2 'd 2));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1288 (.out1(_1220), .in1(_1219), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1271 (.out1(_1203), .in1(_1202), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1235 (.out1(_1167), .in1(_1166), .in2(63 'd 6148914691236517205));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1289 (.out1(_1221), .in1(_1203), .in2(_1220));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1253 (.out1(_1185), .in1(_1184), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1236 (.out1(_1168), .in1(_1159), .in2(_1167));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2862 (.out1(R2863), .clock(clock), .in1(R2862));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3068 (.out1(R3069), .clock(clock), .in1(R3068));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3270 (.out1(R3271), .clock(clock), .in1(R3270));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3517 (.out1(R3518), .clock(clock), .in1(R3517));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3709 (.out1(R3710), .clock(clock), .in1(R3709));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3897 (.out1(R3898), .clock(clock), .in1(R3897));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4130 (.out1(R4131), .clock(clock), .in1(R4130));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4308 (.out1(R4309), .clock(clock), .in1(R4308));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4482 (.out1(R4483), .clock(clock), .in1(R4482));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4701 (.out1(R4702), .clock(clock), .in1(R4701));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4865 (.out1(R4866), .clock(clock), .in1(R4865));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5025 (.out1(R5026), .clock(clock), .in1(R5025));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5230 (.out1(R5231), .clock(clock), .in1(R5230));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5380 (.out1(R5381), .clock(clock), .in1(R5380));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5526 (.out1(R5527), .clock(clock), .in1(R5526));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5717 (.out1(R5718), .clock(clock), .in1(R5717));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5853 (.out1(R5854), .clock(clock), .in1(R5853));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5985 (.out1(R5986), .clock(clock), .in1(R5985));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6161 (.out1(R6162), .clock(clock), .in1(R6161));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6282 (.out1(R6283), .clock(clock), .in1(R6282));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6399 (.out1(R6400), .clock(clock), .in1(R6399));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6562 (.out1(R6563), .clock(clock), .in1(R6562));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6669 (.out1(R6670), .clock(clock), .in1(R6669));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6772 (.out1(R6773), .clock(clock), .in1(R6772));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6920 (.out1(R6921), .clock(clock), .in1(R6920));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7013 (.out1(R7014), .clock(clock), .in1(R7013));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7102 (.out1(R7103), .clock(clock), .in1(R7102));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7236 (.out1(R7237), .clock(clock), .in1(R7236));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7315 (.out1(R7316), .clock(clock), .in1(R7315));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7390 (.out1(R7391), .clock(clock), .in1(R7390));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7510 (.out1(R7511), .clock(clock), .in1(R7510));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7575 (.out1(R7576), .clock(clock), .in1(R7575));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7636 (.out1(R7637), .clock(clock), .in1(R7636));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7742 (.out1(R7743), .clock(clock), .in1(R7742));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7793 (.out1(R7794), .clock(clock), .in1(R7793));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7840 (.out1(R7841), .clock(clock), .in1(R7840));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7932 (.out1(R7933), .clock(clock), .in1(R7932));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7969 (.out1(R7970), .clock(clock), .in1(R7969));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8002 (.out1(R8003), .clock(clock), .in1(R8002));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8080 (.out1(R8081), .clock(clock), .in1(R8080));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8103 (.out1(R8104), .clock(clock), .in1(R8103));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8122 (.out1(R8123), .clock(clock), .in1(R8122));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8177 (.out1(R8178), .clock(clock), .in1(_1151));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8178 (.out1(R8179), .clock(clock), .in1(_1221));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8179 (.out1(R8180), .clock(clock), .in1(_1185));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8180 (.out1(R8181), .clock(clock), .in1(_1168));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1254 (.out1(_1186), .in1(R8180), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1237 (.out1(_1169), .in1(R8181), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op1290 (.out1(_1222), .in1(R8179), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1255 (.out1(_1187), .in1(_1169), .in2(_1186));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1220 (.out1(_1152), .in1(c120_popcnt_2664_D), .in2(R8178));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1291 (.out1(_1223), .in1(_1187), .in2(_1222));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op1292 (.out1(_1224), .in1(_1223), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2863 (.out1(R2864), .clock(clock), .in1(R2863));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3069 (.out1(R3070), .clock(clock), .in1(R3069));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3271 (.out1(R3272), .clock(clock), .in1(R3271));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3518 (.out1(R3519), .clock(clock), .in1(R3518));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3710 (.out1(R3711), .clock(clock), .in1(R3710));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3898 (.out1(R3899), .clock(clock), .in1(R3898));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4131 (.out1(R4132), .clock(clock), .in1(R4131));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4309 (.out1(R4310), .clock(clock), .in1(R4309));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4483 (.out1(R4484), .clock(clock), .in1(R4483));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4702 (.out1(R4703), .clock(clock), .in1(R4702));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4866 (.out1(R4867), .clock(clock), .in1(R4866));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5026 (.out1(R5027), .clock(clock), .in1(R5026));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5231 (.out1(R5232), .clock(clock), .in1(R5231));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5381 (.out1(R5382), .clock(clock), .in1(R5381));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5527 (.out1(R5528), .clock(clock), .in1(R5527));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5718 (.out1(R5719), .clock(clock), .in1(R5718));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5854 (.out1(R5855), .clock(clock), .in1(R5854));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5986 (.out1(R5987), .clock(clock), .in1(R5986));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6162 (.out1(R6163), .clock(clock), .in1(R6162));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6283 (.out1(R6284), .clock(clock), .in1(R6283));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6400 (.out1(R6401), .clock(clock), .in1(R6400));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6563 (.out1(R6564), .clock(clock), .in1(R6563));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6670 (.out1(R6671), .clock(clock), .in1(R6670));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6773 (.out1(R6774), .clock(clock), .in1(R6773));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6921 (.out1(R6922), .clock(clock), .in1(R6921));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7014 (.out1(R7015), .clock(clock), .in1(R7014));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7103 (.out1(R7104), .clock(clock), .in1(R7103));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7237 (.out1(R7238), .clock(clock), .in1(R7237));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7316 (.out1(R7317), .clock(clock), .in1(R7316));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7391 (.out1(R7392), .clock(clock), .in1(R7391));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7511 (.out1(R7512), .clock(clock), .in1(R7511));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7576 (.out1(R7577), .clock(clock), .in1(R7576));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7637 (.out1(R7638), .clock(clock), .in1(R7637));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7743 (.out1(R7744), .clock(clock), .in1(R7743));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7794 (.out1(R7795), .clock(clock), .in1(R7794));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7841 (.out1(R7842), .clock(clock), .in1(R7841));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7933 (.out1(R7934), .clock(clock), .in1(R7933));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7970 (.out1(R7971), .clock(clock), .in1(R7970));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8003 (.out1(R8004), .clock(clock), .in1(R8003));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8081 (.out1(R8082), .clock(clock), .in1(R8081));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8104 (.out1(R8105), .clock(clock), .in1(R8104));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8123 (.out1(R8124), .clock(clock), .in1(R8123));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8181 (.out1(R8182), .clock(clock), .in1(_1152));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8182 (.out1(R8183), .clock(clock), .in1(_1224));
  SRAM op1221 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1153),.ADR(R8182));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op1293 (.out1(_1225), .in1(R8183), .in2(57 'd 72340172838076673));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2864 (.out1(R2865), .clock(clock), .in1(R2864));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3070 (.out1(R3071), .clock(clock), .in1(R3070));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3272 (.out1(R3273), .clock(clock), .in1(R3272));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3519 (.out1(R3520), .clock(clock), .in1(R3519));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3711 (.out1(R3712), .clock(clock), .in1(R3711));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3899 (.out1(R3900), .clock(clock), .in1(R3899));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4132 (.out1(R4133), .clock(clock), .in1(R4132));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4310 (.out1(R4311), .clock(clock), .in1(R4310));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4484 (.out1(R4485), .clock(clock), .in1(R4484));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4703 (.out1(R4704), .clock(clock), .in1(R4703));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4867 (.out1(R4868), .clock(clock), .in1(R4867));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5027 (.out1(R5028), .clock(clock), .in1(R5027));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5232 (.out1(R5233), .clock(clock), .in1(R5232));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5382 (.out1(R5383), .clock(clock), .in1(R5382));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5528 (.out1(R5529), .clock(clock), .in1(R5528));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5719 (.out1(R5720), .clock(clock), .in1(R5719));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5855 (.out1(R5856), .clock(clock), .in1(R5855));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5987 (.out1(R5988), .clock(clock), .in1(R5987));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6163 (.out1(R6164), .clock(clock), .in1(R6163));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6284 (.out1(R6285), .clock(clock), .in1(R6284));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6401 (.out1(R6402), .clock(clock), .in1(R6401));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6564 (.out1(R6565), .clock(clock), .in1(R6564));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6671 (.out1(R6672), .clock(clock), .in1(R6671));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6774 (.out1(R6775), .clock(clock), .in1(R6774));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6922 (.out1(R6923), .clock(clock), .in1(R6922));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7015 (.out1(R7016), .clock(clock), .in1(R7015));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7104 (.out1(R7105), .clock(clock), .in1(R7104));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7238 (.out1(R7239), .clock(clock), .in1(R7238));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7317 (.out1(R7318), .clock(clock), .in1(R7317));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7392 (.out1(R7393), .clock(clock), .in1(R7392));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7512 (.out1(R7513), .clock(clock), .in1(R7512));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7577 (.out1(R7578), .clock(clock), .in1(R7577));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7638 (.out1(R7639), .clock(clock), .in1(R7638));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7744 (.out1(R7745), .clock(clock), .in1(R7744));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7795 (.out1(R7796), .clock(clock), .in1(R7795));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7842 (.out1(R7843), .clock(clock), .in1(R7842));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7934 (.out1(R7935), .clock(clock), .in1(R7934));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7971 (.out1(R7972), .clock(clock), .in1(R7971));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8004 (.out1(R8005), .clock(clock), .in1(R8004));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8082 (.out1(R8083), .clock(clock), .in1(R8082));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8105 (.out1(R8106), .clock(clock), .in1(R8105));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8124 (.out1(R8125), .clock(clock), .in1(R8124));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8183 (.out1(R8184), .clock(clock), .in1(_1153));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8184 (.out1(R8185), .clock(clock), .in1(_1225));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op1294 (.out1(_1226), .in1(R8185), .in2(6 'd 56));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1295 (.out1(_1227), .in1(_1226));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1296 (.out1(ck_idx_2665), .in1(R8184), .in2(_1227));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2865 (.out1(R2866), .clock(clock), .in1(R2865));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3071 (.out1(R3072), .clock(clock), .in1(R3071));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3273 (.out1(R3274), .clock(clock), .in1(R3273));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3520 (.out1(R3521), .clock(clock), .in1(R3520));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3712 (.out1(R3713), .clock(clock), .in1(R3712));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3900 (.out1(R3901), .clock(clock), .in1(R3900));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4133 (.out1(R4134), .clock(clock), .in1(R4133));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4311 (.out1(R4312), .clock(clock), .in1(R4311));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4485 (.out1(R4486), .clock(clock), .in1(R4485));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4704 (.out1(R4705), .clock(clock), .in1(R4704));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4868 (.out1(R4869), .clock(clock), .in1(R4868));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5028 (.out1(R5029), .clock(clock), .in1(R5028));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5233 (.out1(R5234), .clock(clock), .in1(R5233));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5383 (.out1(R5384), .clock(clock), .in1(R5383));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5529 (.out1(R5530), .clock(clock), .in1(R5529));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5720 (.out1(R5721), .clock(clock), .in1(R5720));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5856 (.out1(R5857), .clock(clock), .in1(R5856));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5988 (.out1(R5989), .clock(clock), .in1(R5988));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6164 (.out1(R6165), .clock(clock), .in1(R6164));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6285 (.out1(R6286), .clock(clock), .in1(R6285));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6402 (.out1(R6403), .clock(clock), .in1(R6402));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6565 (.out1(R6566), .clock(clock), .in1(R6565));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6672 (.out1(R6673), .clock(clock), .in1(R6672));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6775 (.out1(R6776), .clock(clock), .in1(R6775));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6923 (.out1(R6924), .clock(clock), .in1(R6923));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7016 (.out1(R7017), .clock(clock), .in1(R7016));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7105 (.out1(R7106), .clock(clock), .in1(R7105));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7239 (.out1(R7240), .clock(clock), .in1(R7239));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7318 (.out1(R7319), .clock(clock), .in1(R7318));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7393 (.out1(R7394), .clock(clock), .in1(R7393));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7513 (.out1(R7514), .clock(clock), .in1(R7513));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7578 (.out1(R7579), .clock(clock), .in1(R7578));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7639 (.out1(R7640), .clock(clock), .in1(R7639));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7745 (.out1(R7746), .clock(clock), .in1(R7745));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7796 (.out1(R7797), .clock(clock), .in1(R7796));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7843 (.out1(R7844), .clock(clock), .in1(R7843));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7935 (.out1(R7936), .clock(clock), .in1(R7935));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7972 (.out1(R7973), .clock(clock), .in1(R7972));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8005 (.out1(R8006), .clock(clock), .in1(R8005));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8083 (.out1(R8084), .clock(clock), .in1(R8083));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8106 (.out1(R8107), .clock(clock), .in1(R8106));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8125 (.out1(R8126), .clock(clock), .in1(R8125));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8185 (.out1(R8186), .clock(clock), .in1(ck_idx_2665));
  LSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(4), .BITSIZE_out1(32), .PRECISION(32)) op1297 (.out1(_1228), .in1(R8186), .in2(4 'd 8));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2866 (.out1(R2867), .clock(clock), .in1(R2866));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3072 (.out1(R3073), .clock(clock), .in1(R3072));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3274 (.out1(R3275), .clock(clock), .in1(R3274));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3521 (.out1(R3522), .clock(clock), .in1(R3521));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3713 (.out1(R3714), .clock(clock), .in1(R3713));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3901 (.out1(R3902), .clock(clock), .in1(R3901));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4134 (.out1(R4135), .clock(clock), .in1(R4134));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4312 (.out1(R4313), .clock(clock), .in1(R4312));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4486 (.out1(R4487), .clock(clock), .in1(R4486));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4705 (.out1(R4706), .clock(clock), .in1(R4705));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4869 (.out1(R4870), .clock(clock), .in1(R4869));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5029 (.out1(R5030), .clock(clock), .in1(R5029));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5234 (.out1(R5235), .clock(clock), .in1(R5234));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5384 (.out1(R5385), .clock(clock), .in1(R5384));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5530 (.out1(R5531), .clock(clock), .in1(R5530));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5721 (.out1(R5722), .clock(clock), .in1(R5721));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5857 (.out1(R5858), .clock(clock), .in1(R5857));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5989 (.out1(R5990), .clock(clock), .in1(R5989));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6165 (.out1(R6166), .clock(clock), .in1(R6165));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6286 (.out1(R6287), .clock(clock), .in1(R6286));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6403 (.out1(R6404), .clock(clock), .in1(R6403));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6566 (.out1(R6567), .clock(clock), .in1(R6566));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6673 (.out1(R6674), .clock(clock), .in1(R6673));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6776 (.out1(R6777), .clock(clock), .in1(R6776));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6924 (.out1(R6925), .clock(clock), .in1(R6924));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7017 (.out1(R7018), .clock(clock), .in1(R7017));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7106 (.out1(R7107), .clock(clock), .in1(R7106));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7240 (.out1(R7241), .clock(clock), .in1(R7240));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7319 (.out1(R7320), .clock(clock), .in1(R7319));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7394 (.out1(R7395), .clock(clock), .in1(R7394));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7514 (.out1(R7515), .clock(clock), .in1(R7514));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7579 (.out1(R7580), .clock(clock), .in1(R7579));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7640 (.out1(R7641), .clock(clock), .in1(R7640));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7746 (.out1(R7747), .clock(clock), .in1(R7746));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7797 (.out1(R7798), .clock(clock), .in1(R7797));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7844 (.out1(R7845), .clock(clock), .in1(R7844));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7936 (.out1(R7937), .clock(clock), .in1(R7936));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7973 (.out1(R7974), .clock(clock), .in1(R7973));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8006 (.out1(R8007), .clock(clock), .in1(R8006));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8084 (.out1(R8085), .clock(clock), .in1(R8084));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8107 (.out1(R8108), .clock(clock), .in1(R8107));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8126 (.out1(R8127), .clock(clock), .in1(R8126));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8186 (.out1(R8187), .clock(clock), .in1(_1228));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1298 (.out1(_1229), .in1(ip2_2595_D));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(8), .BITSIZE_out1(32)) op1299 (.out1(_1230), .in1(_1229), .in2(8 'd 255));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1300 (.out1(idx_sail_2666), .in1(R8187), .in2(_1230));
  RSHIFT_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(3), .BITSIZE_out1(32), .PRECISION(32)) op1301 (.out1(idx_2667), .in1(idx_sail_2666), .in2(3 'd 6));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2867 (.out1(R2868), .clock(clock), .in1(R2867));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3073 (.out1(R3074), .clock(clock), .in1(R3073));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3275 (.out1(R3276), .clock(clock), .in1(R3275));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3522 (.out1(R3523), .clock(clock), .in1(R3522));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3714 (.out1(R3715), .clock(clock), .in1(R3714));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3902 (.out1(R3903), .clock(clock), .in1(R3902));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4135 (.out1(R4136), .clock(clock), .in1(R4135));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4313 (.out1(R4314), .clock(clock), .in1(R4313));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4487 (.out1(R4488), .clock(clock), .in1(R4487));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4706 (.out1(R4707), .clock(clock), .in1(R4706));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4870 (.out1(R4871), .clock(clock), .in1(R4870));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5030 (.out1(R5031), .clock(clock), .in1(R5030));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5235 (.out1(R5236), .clock(clock), .in1(R5235));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5385 (.out1(R5386), .clock(clock), .in1(R5385));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5531 (.out1(R5532), .clock(clock), .in1(R5531));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5722 (.out1(R5723), .clock(clock), .in1(R5722));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5858 (.out1(R5859), .clock(clock), .in1(R5858));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5990 (.out1(R5991), .clock(clock), .in1(R5990));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6166 (.out1(R6167), .clock(clock), .in1(R6166));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6287 (.out1(R6288), .clock(clock), .in1(R6287));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6404 (.out1(R6405), .clock(clock), .in1(R6404));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6567 (.out1(R6568), .clock(clock), .in1(R6567));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6674 (.out1(R6675), .clock(clock), .in1(R6674));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6777 (.out1(R6778), .clock(clock), .in1(R6777));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6925 (.out1(R6926), .clock(clock), .in1(R6925));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7018 (.out1(R7019), .clock(clock), .in1(R7018));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7107 (.out1(R7108), .clock(clock), .in1(R7107));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7241 (.out1(R7242), .clock(clock), .in1(R7241));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7320 (.out1(R7321), .clock(clock), .in1(R7320));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7395 (.out1(R7396), .clock(clock), .in1(R7395));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7515 (.out1(R7516), .clock(clock), .in1(R7515));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7580 (.out1(R7581), .clock(clock), .in1(R7580));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7641 (.out1(R7642), .clock(clock), .in1(R7641));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7747 (.out1(R7748), .clock(clock), .in1(R7747));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7798 (.out1(R7799), .clock(clock), .in1(R7798));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7845 (.out1(R7846), .clock(clock), .in1(R7845));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7937 (.out1(R7938), .clock(clock), .in1(R7937));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7974 (.out1(R7975), .clock(clock), .in1(R7974));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8007 (.out1(R8008), .clock(clock), .in1(R8007));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8085 (.out1(R8086), .clock(clock), .in1(R8085));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8108 (.out1(R8109), .clock(clock), .in1(R8108));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8127 (.out1(R8128), .clock(clock), .in1(R8127));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8187 (.out1(R8188), .clock(clock), .in1(idx_sail_2666));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8190 (.out1(R8191), .clock(clock), .in1(idx_2667));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2015 (.out1(_1919), .in1(R6167));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1926 (.out1(_1833), .in1(R6568));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1837 (.out1(_1747), .in1(R6926));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1748 (.out1(_1661), .in1(R7242));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1659 (.out1(_1575), .in1(R7516));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1570 (.out1(_1489), .in1(R7748));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1481 (.out1(_1403), .in1(R7938));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1392 (.out1(_1317), .in1(R8086));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1303 (.out1(_1231), .in1(R8191));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2016 (.out1(_1920), .in1(_1919), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1927 (.out1(_1834), .in1(_1833), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1838 (.out1(_1748), .in1(_1747), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1749 (.out1(_1662), .in1(_1661), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1660 (.out1(_1576), .in1(_1575), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1571 (.out1(_1490), .in1(_1489), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1482 (.out1(_1404), .in1(_1403), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1393 (.out1(_1318), .in1(_1317), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1304 (.out1(_1232), .in1(_1231), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2868 (.out1(R2869), .clock(clock), .in1(R2868));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3074 (.out1(R3075), .clock(clock), .in1(R3074));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3276 (.out1(R3277), .clock(clock), .in1(R3276));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3523 (.out1(R3524), .clock(clock), .in1(R3523));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3715 (.out1(R3716), .clock(clock), .in1(R3715));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3903 (.out1(R3904), .clock(clock), .in1(R3903));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4136 (.out1(R4137), .clock(clock), .in1(R4136));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4314 (.out1(R4315), .clock(clock), .in1(R4314));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4488 (.out1(R4489), .clock(clock), .in1(R4488));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4707 (.out1(R4708), .clock(clock), .in1(R4707));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4871 (.out1(R4872), .clock(clock), .in1(R4871));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5031 (.out1(R5032), .clock(clock), .in1(R5031));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5236 (.out1(R5237), .clock(clock), .in1(R5236));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5386 (.out1(R5387), .clock(clock), .in1(R5386));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5532 (.out1(R5533), .clock(clock), .in1(R5532));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5723 (.out1(R5724), .clock(clock), .in1(R5723));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5859 (.out1(R5860), .clock(clock), .in1(R5859));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5991 (.out1(R5992), .clock(clock), .in1(R5991));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6167 (.out1(R6168), .clock(clock), .in1(R6167));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6288 (.out1(R6289), .clock(clock), .in1(R6288));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6405 (.out1(R6406), .clock(clock), .in1(R6405));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6568 (.out1(R6569), .clock(clock), .in1(R6568));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6675 (.out1(R6676), .clock(clock), .in1(R6675));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6778 (.out1(R6779), .clock(clock), .in1(R6778));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6926 (.out1(R6927), .clock(clock), .in1(R6926));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7019 (.out1(R7020), .clock(clock), .in1(R7019));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7108 (.out1(R7109), .clock(clock), .in1(R7108));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7242 (.out1(R7243), .clock(clock), .in1(R7242));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7321 (.out1(R7322), .clock(clock), .in1(R7321));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7396 (.out1(R7397), .clock(clock), .in1(R7396));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7516 (.out1(R7517), .clock(clock), .in1(R7516));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7581 (.out1(R7582), .clock(clock), .in1(R7581));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7642 (.out1(R7643), .clock(clock), .in1(R7642));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7748 (.out1(R7749), .clock(clock), .in1(R7748));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7799 (.out1(R7800), .clock(clock), .in1(R7799));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7846 (.out1(R7847), .clock(clock), .in1(R7846));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7938 (.out1(R7939), .clock(clock), .in1(R7938));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7975 (.out1(R7976), .clock(clock), .in1(R7975));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8008 (.out1(R8009), .clock(clock), .in1(R8008));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8086 (.out1(R8087), .clock(clock), .in1(R8086));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8109 (.out1(R8110), .clock(clock), .in1(R8109));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8128 (.out1(R8129), .clock(clock), .in1(R8128));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8188 (.out1(R8189), .clock(clock), .in1(R8188));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8191 (.out1(R8192), .clock(clock), .in1(R8191));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8199 (.out1(R8200), .clock(clock), .in1(_1920));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8200 (.out1(R8201), .clock(clock), .in1(_1834));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8201 (.out1(R8202), .clock(clock), .in1(_1748));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8202 (.out1(R8203), .clock(clock), .in1(_1662));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8203 (.out1(R8204), .clock(clock), .in1(_1576));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8204 (.out1(R8205), .clock(clock), .in1(_1490));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8205 (.out1(R8206), .clock(clock), .in1(_1404));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8206 (.out1(R8207), .clock(clock), .in1(_1318));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8207 (.out1(R8208), .clock(clock), .in1(_1232));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2549 (.out1(_2435), .in1(R2869));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2460 (.out1(_2349), .in1(R3524));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2371 (.out1(_2263), .in1(R4137));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2282 (.out1(_2177), .in1(R4708));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2193 (.out1(_2091), .in1(R5237));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2104 (.out1(_2005), .in1(R5724));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2550 (.out1(_2436), .in1(_2435), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2461 (.out1(_2350), .in1(_2349), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2372 (.out1(_2264), .in1(_2263), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2283 (.out1(_2178), .in1(_2177), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2194 (.out1(_2092), .in1(_2091), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2105 (.out1(_2006), .in1(_2005), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2017 (.out1(_1921), .in1(b64_bitmap_2589_D), .in2(R8200));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1928 (.out1(_1835), .in1(b72_bitmap_2600_D), .in2(R8201));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1839 (.out1(_1749), .in1(b80_bitmap_2610_D), .in2(R8202));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1750 (.out1(_1663), .in1(b88_bitmap_2620_D), .in2(R8203));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1661 (.out1(_1577), .in1(b96_bitmap_2630_D), .in2(R8204));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1572 (.out1(_1491), .in1(b104_bitmap_2640_D), .in2(R8205));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1483 (.out1(_1405), .in1(b112_bitmap_2650_D), .in2(R8206));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1394 (.out1(_1319), .in1(b120_bitmap_2660_D), .in2(R8207));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1305 (.out1(_1233), .in1(b128_bitmap_2669_D), .in2(R8208));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2869 (.out1(R2870), .clock(clock), .in1(R2869));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3075 (.out1(R3076), .clock(clock), .in1(R3075));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3277 (.out1(R3278), .clock(clock), .in1(R3277));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3524 (.out1(R3525), .clock(clock), .in1(R3524));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3716 (.out1(R3717), .clock(clock), .in1(R3716));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3904 (.out1(R3905), .clock(clock), .in1(R3904));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4137 (.out1(R4138), .clock(clock), .in1(R4137));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4315 (.out1(R4316), .clock(clock), .in1(R4315));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4489 (.out1(R4490), .clock(clock), .in1(R4489));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4708 (.out1(R4709), .clock(clock), .in1(R4708));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4872 (.out1(R4873), .clock(clock), .in1(R4872));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5032 (.out1(R5033), .clock(clock), .in1(R5032));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5237 (.out1(R5238), .clock(clock), .in1(R5237));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5387 (.out1(R5388), .clock(clock), .in1(R5387));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5533 (.out1(R5534), .clock(clock), .in1(R5533));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5724 (.out1(R5725), .clock(clock), .in1(R5724));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5860 (.out1(R5861), .clock(clock), .in1(R5860));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5992 (.out1(R5993), .clock(clock), .in1(R5992));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6168 (.out1(R6169), .clock(clock), .in1(R6168));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6289 (.out1(R6290), .clock(clock), .in1(R6289));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6406 (.out1(R6407), .clock(clock), .in1(R6406));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6569 (.out1(R6570), .clock(clock), .in1(R6569));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6676 (.out1(R6677), .clock(clock), .in1(R6676));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6779 (.out1(R6780), .clock(clock), .in1(R6779));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6927 (.out1(R6928), .clock(clock), .in1(R6927));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7020 (.out1(R7021), .clock(clock), .in1(R7020));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7109 (.out1(R7110), .clock(clock), .in1(R7109));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7243 (.out1(R7244), .clock(clock), .in1(R7243));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7322 (.out1(R7323), .clock(clock), .in1(R7322));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7397 (.out1(R7398), .clock(clock), .in1(R7397));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7517 (.out1(R7518), .clock(clock), .in1(R7517));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7582 (.out1(R7583), .clock(clock), .in1(R7582));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7643 (.out1(R7644), .clock(clock), .in1(R7643));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7749 (.out1(R7750), .clock(clock), .in1(R7749));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7800 (.out1(R7801), .clock(clock), .in1(R7800));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7847 (.out1(R7848), .clock(clock), .in1(R7847));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7939 (.out1(R7940), .clock(clock), .in1(R7939));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7976 (.out1(R7977), .clock(clock), .in1(R7976));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8009 (.out1(R8010), .clock(clock), .in1(R8009));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8087 (.out1(R8088), .clock(clock), .in1(R8087));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8110 (.out1(R8111), .clock(clock), .in1(R8110));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8129 (.out1(R8130), .clock(clock), .in1(R8129));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8189 (.out1(R8190), .clock(clock), .in1(R8189));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8192 (.out1(R8193), .clock(clock), .in1(R8192));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8208 (.out1(R8209), .clock(clock), .in1(_2436));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8209 (.out1(R8210), .clock(clock), .in1(_2350));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8210 (.out1(R8211), .clock(clock), .in1(_2264));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8211 (.out1(R8212), .clock(clock), .in1(_2178));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8212 (.out1(R8213), .clock(clock), .in1(_2092));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8213 (.out1(R8214), .clock(clock), .in1(_2006));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8214 (.out1(R8215), .clock(clock), .in1(_1921));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8215 (.out1(R8216), .clock(clock), .in1(_1835));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8216 (.out1(R8217), .clock(clock), .in1(_1749));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8217 (.out1(R8218), .clock(clock), .in1(_1663));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8218 (.out1(R8219), .clock(clock), .in1(_1577));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8219 (.out1(R8220), .clock(clock), .in1(_1491));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8220 (.out1(R8221), .clock(clock), .in1(_1405));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8221 (.out1(R8222), .clock(clock), .in1(_1319));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8222 (.out1(R8223), .clock(clock), .in1(_1233));
  SRAM op2018 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1922),.ADR(R8215));
  SRAM op1929 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1836),.ADR(R8216));
  SRAM op1840 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1750),.ADR(R8217));
  SRAM op1751 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1664),.ADR(R8218));
  SRAM op1662 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1578),.ADR(R8219));
  SRAM op1573 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1492),.ADR(R8220));
  SRAM op1484 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1406),.ADR(R8221));
  SRAM op1395 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1320),.ADR(R8222));
  SRAM op1306 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1234),.ADR(R8223));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2551 (.out1(_2437), .in1(b16_bitmap_2528_D), .in2(R8209));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2462 (.out1(_2351), .in1(b24_bitmap_2539_D), .in2(R8210));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2373 (.out1(_2265), .in1(b32_bitmap_2549_D), .in2(R8211));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2284 (.out1(_2179), .in1(b40_bitmap_2559_D), .in2(R8212));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2195 (.out1(_2093), .in1(b48_bitmap_2569_D), .in2(R8213));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2106 (.out1(_2007), .in1(b56_bitmap_2579_D), .in2(R8214));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op1302 (.out1(off_2668), .in1(R8190), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2019 (.out1(_1923), .in1(64 'd 9223372036854775808), .in2(R6290));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1930 (.out1(_1837), .in1(64 'd 9223372036854775808), .in2(R6677));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1841 (.out1(_1751), .in1(64 'd 9223372036854775808), .in2(R7021));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1752 (.out1(_1665), .in1(64 'd 9223372036854775808), .in2(R7323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1663 (.out1(_1579), .in1(64 'd 9223372036854775808), .in2(R7583));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1574 (.out1(_1493), .in1(64 'd 9223372036854775808), .in2(R7801));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1485 (.out1(_1407), .in1(64 'd 9223372036854775808), .in2(R7977));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1396 (.out1(_1321), .in1(64 'd 9223372036854775808), .in2(R8111));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1307 (.out1(_1235), .in1(64 'd 9223372036854775808), .in2(off_2668));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2870 (.out1(R2871), .clock(clock), .in1(R2870));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3076 (.out1(R3077), .clock(clock), .in1(R3076));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3278 (.out1(R3279), .clock(clock), .in1(R3278));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3525 (.out1(R3526), .clock(clock), .in1(R3525));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3717 (.out1(R3718), .clock(clock), .in1(R3717));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3905 (.out1(R3906), .clock(clock), .in1(R3905));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4138 (.out1(R4139), .clock(clock), .in1(R4138));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4316 (.out1(R4317), .clock(clock), .in1(R4316));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4490 (.out1(R4491), .clock(clock), .in1(R4490));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4709 (.out1(R4710), .clock(clock), .in1(R4709));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4873 (.out1(R4874), .clock(clock), .in1(R4873));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5033 (.out1(R5034), .clock(clock), .in1(R5033));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5238 (.out1(R5239), .clock(clock), .in1(R5238));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5388 (.out1(R5389), .clock(clock), .in1(R5388));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5534 (.out1(R5535), .clock(clock), .in1(R5534));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5725 (.out1(R5726), .clock(clock), .in1(R5725));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5861 (.out1(R5862), .clock(clock), .in1(R5861));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5993 (.out1(R5994), .clock(clock), .in1(R5993));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6169 (.out1(R6170), .clock(clock), .in1(R6169));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6290 (.out1(R6291), .clock(clock), .in1(R6290));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6407 (.out1(R6408), .clock(clock), .in1(R6407));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6570 (.out1(R6571), .clock(clock), .in1(R6570));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6677 (.out1(R6678), .clock(clock), .in1(R6677));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6780 (.out1(R6781), .clock(clock), .in1(R6780));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6928 (.out1(R6929), .clock(clock), .in1(R6928));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7021 (.out1(R7022), .clock(clock), .in1(R7021));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7110 (.out1(R7111), .clock(clock), .in1(R7110));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7244 (.out1(R7245), .clock(clock), .in1(R7244));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7323 (.out1(R7324), .clock(clock), .in1(R7323));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7398 (.out1(R7399), .clock(clock), .in1(R7398));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7518 (.out1(R7519), .clock(clock), .in1(R7518));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7583 (.out1(R7584), .clock(clock), .in1(R7583));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7644 (.out1(R7645), .clock(clock), .in1(R7644));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7750 (.out1(R7751), .clock(clock), .in1(R7750));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7801 (.out1(R7802), .clock(clock), .in1(R7801));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7848 (.out1(R7849), .clock(clock), .in1(R7848));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7940 (.out1(R7941), .clock(clock), .in1(R7940));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7977 (.out1(R7978), .clock(clock), .in1(R7977));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8010 (.out1(R8011), .clock(clock), .in1(R8010));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8088 (.out1(R8089), .clock(clock), .in1(R8088));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8111 (.out1(R8112), .clock(clock), .in1(R8111));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8130 (.out1(R8131), .clock(clock), .in1(R8130));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8193 (.out1(R8194), .clock(clock), .in1(R8193));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8223 (.out1(R8224), .clock(clock), .in1(_1922));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8224 (.out1(R8225), .clock(clock), .in1(_1836));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8225 (.out1(R8226), .clock(clock), .in1(_1750));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8226 (.out1(R8227), .clock(clock), .in1(_1664));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8227 (.out1(R8228), .clock(clock), .in1(_1578));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8228 (.out1(R8229), .clock(clock), .in1(_1492));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8229 (.out1(R8230), .clock(clock), .in1(_1406));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8230 (.out1(R8231), .clock(clock), .in1(_1320));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8231 (.out1(R8232), .clock(clock), .in1(_1234));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8232 (.out1(R8233), .clock(clock), .in1(_2437));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8233 (.out1(R8234), .clock(clock), .in1(_2351));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8234 (.out1(R8235), .clock(clock), .in1(_2265));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8235 (.out1(R8236), .clock(clock), .in1(_2179));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8236 (.out1(R8237), .clock(clock), .in1(_2093));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8237 (.out1(R8238), .clock(clock), .in1(_2007));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8238 (.out1(R8239), .clock(clock), .in1(off_2668));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8243 (.out1(R8244), .clock(clock), .in1(_1923));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8244 (.out1(R8245), .clock(clock), .in1(_1837));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8245 (.out1(R8246), .clock(clock), .in1(_1751));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8246 (.out1(R8247), .clock(clock), .in1(_1665));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8247 (.out1(R8248), .clock(clock), .in1(_1579));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8248 (.out1(R8249), .clock(clock), .in1(_1493));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8249 (.out1(R8250), .clock(clock), .in1(_1407));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8250 (.out1(R8251), .clock(clock), .in1(_1321));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8251 (.out1(R8252), .clock(clock), .in1(_1235));
  SRAM op2552 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2438),.ADR(R8233));
  SRAM op2463 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2352),.ADR(R8234));
  SRAM op2374 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2266),.ADR(R8235));
  SRAM op2285 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2180),.ADR(R8236));
  SRAM op2196 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2094),.ADR(R8237));
  SRAM op2107 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2008),.ADR(R8238));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2020 (.out1(_1924), .in1(R8224), .in2(R8244));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1931 (.out1(_1838), .in1(R8225), .in2(R8245));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1842 (.out1(_1752), .in1(R8226), .in2(R8246));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1753 (.out1(_1666), .in1(R8227), .in2(R8247));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1664 (.out1(_1580), .in1(R8228), .in2(R8248));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1575 (.out1(_1494), .in1(R8229), .in2(R8249));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1486 (.out1(_1408), .in1(R8230), .in2(R8250));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1397 (.out1(_1322), .in1(R8231), .in2(R8251));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1308 (.out1(_1236), .in1(R8232), .in2(R8252));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op2021 (.out1(ifout2021), .in1(_1924), .in2(1 'd 0));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op1932 (.out1(ifout1932), .in1(_1838), .in2(1 'd 0));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op1843 (.out1(ifout1843), .in1(_1752), .in2(1 'd 0));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op1754 (.out1(ifout1754), .in1(_1666), .in2(1 'd 0));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op1665 (.out1(ifout1665), .in1(_1580), .in2(1 'd 0));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op1576 (.out1(ifout1576), .in1(_1494), .in2(1 'd 0));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op1487 (.out1(ifout1487), .in1(_1408), .in2(1 'd 0));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op1398 (.out1(ifout1398), .in1(_1322), .in2(1 'd 0));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op1309 (.out1(ifout1309), .in1(_1236), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2082 (.out1(_1985), .in1(R6170));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1993 (.out1(_1899), .in1(R6571));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1904 (.out1(_1813), .in1(R6929));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1815 (.out1(_1727), .in1(R7245));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1726 (.out1(_1641), .in1(R7519));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1637 (.out1(_1555), .in1(R7751));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1548 (.out1(_1469), .in1(R7941));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1459 (.out1(_1383), .in1(R8089));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1370 (.out1(_1297), .in1(R8194));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2083 (.out1(_1986), .in1(_1985), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1994 (.out1(_1900), .in1(_1899), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1905 (.out1(_1814), .in1(_1813), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1816 (.out1(_1728), .in1(_1727), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1727 (.out1(_1642), .in1(_1641), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1638 (.out1(_1556), .in1(_1555), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1549 (.out1(_1470), .in1(_1469), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1460 (.out1(_1384), .in1(_1383), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1371 (.out1(_1298), .in1(_1297), .in2(2 'd 3));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2553 (.out1(_2439), .in1(64 'd 9223372036854775808), .in2(R3077));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2464 (.out1(_2353), .in1(64 'd 9223372036854775808), .in2(R3718));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2375 (.out1(_2267), .in1(64 'd 9223372036854775808), .in2(R4317));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2286 (.out1(_2181), .in1(64 'd 9223372036854775808), .in2(R4874));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2197 (.out1(_2095), .in1(64 'd 9223372036854775808), .in2(R5389));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2108 (.out1(_2009), .in1(64 'd 9223372036854775808), .in2(R5862));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2871 (.out1(R2872), .clock(clock), .in1(R2871));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3077 (.out1(R3078), .clock(clock), .in1(R3077));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3279 (.out1(R3280), .clock(clock), .in1(R3279));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3526 (.out1(R3527), .clock(clock), .in1(R3526));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3718 (.out1(R3719), .clock(clock), .in1(R3718));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3906 (.out1(R3907), .clock(clock), .in1(R3906));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4139 (.out1(R4140), .clock(clock), .in1(R4139));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4317 (.out1(R4318), .clock(clock), .in1(R4317));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4491 (.out1(R4492), .clock(clock), .in1(R4491));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4710 (.out1(R4711), .clock(clock), .in1(R4710));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4874 (.out1(R4875), .clock(clock), .in1(R4874));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5034 (.out1(R5035), .clock(clock), .in1(R5034));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5239 (.out1(R5240), .clock(clock), .in1(R5239));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5389 (.out1(R5390), .clock(clock), .in1(R5389));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5535 (.out1(R5536), .clock(clock), .in1(R5535));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5726 (.out1(R5727), .clock(clock), .in1(R5726));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5862 (.out1(R5863), .clock(clock), .in1(R5862));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5994 (.out1(R5995), .clock(clock), .in1(R5994));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6170 (.out1(R6171), .clock(clock), .in1(R6170));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6291 (.out1(R6292), .clock(clock), .in1(R6291));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6408 (.out1(R6409), .clock(clock), .in1(R6408));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6571 (.out1(R6572), .clock(clock), .in1(R6571));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6678 (.out1(R6679), .clock(clock), .in1(R6678));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6781 (.out1(R6782), .clock(clock), .in1(R6781));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6929 (.out1(R6930), .clock(clock), .in1(R6929));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7022 (.out1(R7023), .clock(clock), .in1(R7022));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7111 (.out1(R7112), .clock(clock), .in1(R7111));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7245 (.out1(R7246), .clock(clock), .in1(R7245));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7324 (.out1(R7325), .clock(clock), .in1(R7324));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7399 (.out1(R7400), .clock(clock), .in1(R7399));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7519 (.out1(R7520), .clock(clock), .in1(R7519));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7584 (.out1(R7585), .clock(clock), .in1(R7584));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7645 (.out1(R7646), .clock(clock), .in1(R7645));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7751 (.out1(R7752), .clock(clock), .in1(R7751));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7802 (.out1(R7803), .clock(clock), .in1(R7802));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7849 (.out1(R7850), .clock(clock), .in1(R7849));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7941 (.out1(R7942), .clock(clock), .in1(R7941));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7978 (.out1(R7979), .clock(clock), .in1(R7978));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8011 (.out1(R8012), .clock(clock), .in1(R8011));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8089 (.out1(R8090), .clock(clock), .in1(R8089));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8112 (.out1(R8113), .clock(clock), .in1(R8112));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8131 (.out1(R8132), .clock(clock), .in1(R8131));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8194 (.out1(R8195), .clock(clock), .in1(R8194));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8239 (.out1(R8240), .clock(clock), .in1(R8239));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8252 (.out1(R8253), .clock(clock), .in1(_2438));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8253 (.out1(R8254), .clock(clock), .in1(_2352));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8254 (.out1(R8255), .clock(clock), .in1(_2266));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8255 (.out1(R8256), .clock(clock), .in1(_2180));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8256 (.out1(R8257), .clock(clock), .in1(_2094));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8257 (.out1(R8258), .clock(clock), .in1(_2008));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8258 (.out1(R8259), .clock(clock), .in1(ifout2021));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8269 (.out1(R8270), .clock(clock), .in1(ifout1932));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8280 (.out1(R8281), .clock(clock), .in1(ifout1843));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8291 (.out1(R8292), .clock(clock), .in1(ifout1754));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8302 (.out1(R8303), .clock(clock), .in1(ifout1665));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8313 (.out1(R8314), .clock(clock), .in1(ifout1576));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8324 (.out1(R8325), .clock(clock), .in1(ifout1487));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8335 (.out1(R8336), .clock(clock), .in1(ifout1398));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8346 (.out1(R8347), .clock(clock), .in1(ifout1309));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8357 (.out1(R8358), .clock(clock), .in1(_1986));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8358 (.out1(R8359), .clock(clock), .in1(_1900));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8359 (.out1(R8360), .clock(clock), .in1(_1814));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8360 (.out1(R8361), .clock(clock), .in1(_1728));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8361 (.out1(R8362), .clock(clock), .in1(_1642));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8362 (.out1(R8363), .clock(clock), .in1(_1556));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8363 (.out1(R8364), .clock(clock), .in1(_1470));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8364 (.out1(R8365), .clock(clock), .in1(_1384));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8365 (.out1(R8366), .clock(clock), .in1(_1298));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8366 (.out1(R8367), .clock(clock), .in1(_2439));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8367 (.out1(R8368), .clock(clock), .in1(_2353));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8368 (.out1(R8369), .clock(clock), .in1(_2267));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8369 (.out1(R8370), .clock(clock), .in1(_2181));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8370 (.out1(R8371), .clock(clock), .in1(_2095));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8371 (.out1(R8372), .clock(clock), .in1(_2009));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2554 (.out1(_2440), .in1(R8253), .in2(R8367));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2465 (.out1(_2354), .in1(R8254), .in2(R8368));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2376 (.out1(_2268), .in1(R8255), .in2(R8369));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2287 (.out1(_2182), .in1(R8256), .in2(R8370));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2198 (.out1(_2096), .in1(R8257), .in2(R8371));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2109 (.out1(_2010), .in1(R8258), .in2(R8372));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op2555 (.out1(ifout2555), .in1(_2440), .in2(1 'd 0));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op2466 (.out1(ifout2466), .in1(_2354), .in2(1 'd 0));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op2377 (.out1(ifout2377), .in1(_2268), .in2(1 'd 0));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op2288 (.out1(ifout2288), .in1(_2182), .in2(1 'd 0));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op2199 (.out1(ifout2199), .in1(_2096), .in2(1 'd 0));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op2110 (.out1(ifout2110), .in1(_2010), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2616 (.out1(_2501), .in1(R2872));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2527 (.out1(_2415), .in1(R3527));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2438 (.out1(_2329), .in1(R4140));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2349 (.out1(_2243), .in1(R4711));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2260 (.out1(_2157), .in1(R5240));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2171 (.out1(_2071), .in1(R5727));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2076 (.out1(_1979), .in1(R6171));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2066 (.out1(_1969), .in1(R6171));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2060 (.out1(_1963), .in1(R6171));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2048 (.out1(_1951), .in1(R6171));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2042 (.out1(_1945), .in1(R6171));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2032 (.out1(_1935), .in1(R6171));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1987 (.out1(_1893), .in1(R6572));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1977 (.out1(_1883), .in1(R6572));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1971 (.out1(_1877), .in1(R6572));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1959 (.out1(_1865), .in1(R6572));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1953 (.out1(_1859), .in1(R6572));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1943 (.out1(_1849), .in1(R6572));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1898 (.out1(_1807), .in1(R6930));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1888 (.out1(_1797), .in1(R6930));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1882 (.out1(_1791), .in1(R6930));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1870 (.out1(_1779), .in1(R6930));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1864 (.out1(_1773), .in1(R6930));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1854 (.out1(_1763), .in1(R6930));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1809 (.out1(_1721), .in1(R7246));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1799 (.out1(_1711), .in1(R7246));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1793 (.out1(_1705), .in1(R7246));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1781 (.out1(_1693), .in1(R7246));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1775 (.out1(_1687), .in1(R7246));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1765 (.out1(_1677), .in1(R7246));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1720 (.out1(_1635), .in1(R7520));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1710 (.out1(_1625), .in1(R7520));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1704 (.out1(_1619), .in1(R7520));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1692 (.out1(_1607), .in1(R7520));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1686 (.out1(_1601), .in1(R7520));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1676 (.out1(_1591), .in1(R7520));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1631 (.out1(_1549), .in1(R7752));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1621 (.out1(_1539), .in1(R7752));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1615 (.out1(_1533), .in1(R7752));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1603 (.out1(_1521), .in1(R7752));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1597 (.out1(_1515), .in1(R7752));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1587 (.out1(_1505), .in1(R7752));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1542 (.out1(_1463), .in1(R7942));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1532 (.out1(_1453), .in1(R7942));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1526 (.out1(_1447), .in1(R7942));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1514 (.out1(_1435), .in1(R7942));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1508 (.out1(_1429), .in1(R7942));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1498 (.out1(_1419), .in1(R7942));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1453 (.out1(_1377), .in1(R8090));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1443 (.out1(_1367), .in1(R8090));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1437 (.out1(_1361), .in1(R8090));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1425 (.out1(_1349), .in1(R8090));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1419 (.out1(_1343), .in1(R8090));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1409 (.out1(_1333), .in1(R8090));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1364 (.out1(_1291), .in1(R8195));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1354 (.out1(_1281), .in1(R8195));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1348 (.out1(_1275), .in1(R8195));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1336 (.out1(_1263), .in1(R8195));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1330 (.out1(_1257), .in1(R8195));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1320 (.out1(_1247), .in1(R8195));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2617 (.out1(_2502), .in1(_2501), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2528 (.out1(_2416), .in1(_2415), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2439 (.out1(_2330), .in1(_2329), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2350 (.out1(_2244), .in1(_2243), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2261 (.out1(_2158), .in1(_2157), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2172 (.out1(_2072), .in1(_2071), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2077 (.out1(_1980), .in1(_1979), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2067 (.out1(_1970), .in1(_1969), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2061 (.out1(_1964), .in1(_1963), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2049 (.out1(_1952), .in1(_1951), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2043 (.out1(_1946), .in1(_1945), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2033 (.out1(_1936), .in1(_1935), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1988 (.out1(_1894), .in1(_1893), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1978 (.out1(_1884), .in1(_1883), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1972 (.out1(_1878), .in1(_1877), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1960 (.out1(_1866), .in1(_1865), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1954 (.out1(_1860), .in1(_1859), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1944 (.out1(_1850), .in1(_1849), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1899 (.out1(_1808), .in1(_1807), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1889 (.out1(_1798), .in1(_1797), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1883 (.out1(_1792), .in1(_1791), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1871 (.out1(_1780), .in1(_1779), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1865 (.out1(_1774), .in1(_1773), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1855 (.out1(_1764), .in1(_1763), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1810 (.out1(_1722), .in1(_1721), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1800 (.out1(_1712), .in1(_1711), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1794 (.out1(_1706), .in1(_1705), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1782 (.out1(_1694), .in1(_1693), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1776 (.out1(_1688), .in1(_1687), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1766 (.out1(_1678), .in1(_1677), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1721 (.out1(_1636), .in1(_1635), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1711 (.out1(_1626), .in1(_1625), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1705 (.out1(_1620), .in1(_1619), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1693 (.out1(_1608), .in1(_1607), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1687 (.out1(_1602), .in1(_1601), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1677 (.out1(_1592), .in1(_1591), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1632 (.out1(_1550), .in1(_1549), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1622 (.out1(_1540), .in1(_1539), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1616 (.out1(_1534), .in1(_1533), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1604 (.out1(_1522), .in1(_1521), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1598 (.out1(_1516), .in1(_1515), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1588 (.out1(_1506), .in1(_1505), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1543 (.out1(_1464), .in1(_1463), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1533 (.out1(_1454), .in1(_1453), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1527 (.out1(_1448), .in1(_1447), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1515 (.out1(_1436), .in1(_1435), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1509 (.out1(_1430), .in1(_1429), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1499 (.out1(_1420), .in1(_1419), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1454 (.out1(_1378), .in1(_1377), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1444 (.out1(_1368), .in1(_1367), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1438 (.out1(_1362), .in1(_1361), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1426 (.out1(_1350), .in1(_1349), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1420 (.out1(_1344), .in1(_1343), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1410 (.out1(_1334), .in1(_1333), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1365 (.out1(_1292), .in1(_1291), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1355 (.out1(_1282), .in1(_1281), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1349 (.out1(_1276), .in1(_1275), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1337 (.out1(_1264), .in1(_1263), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1331 (.out1(_1258), .in1(_1257), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1321 (.out1(_1248), .in1(_1247), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2084 (.out1(_1987), .in1(b64_bitmap_2589_D), .in2(R8358));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1995 (.out1(_1901), .in1(b72_bitmap_2600_D), .in2(R8359));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1906 (.out1(_1815), .in1(b80_bitmap_2610_D), .in2(R8360));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1817 (.out1(_1729), .in1(b88_bitmap_2620_D), .in2(R8361));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1728 (.out1(_1643), .in1(b96_bitmap_2630_D), .in2(R8362));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1639 (.out1(_1557), .in1(b104_bitmap_2640_D), .in2(R8363));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1550 (.out1(_1471), .in1(b112_bitmap_2650_D), .in2(R8364));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1461 (.out1(_1385), .in1(b120_bitmap_2660_D), .in2(R8365));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1372 (.out1(_1299), .in1(b128_bitmap_2669_D), .in2(R8366));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2872 (.out1(R2873), .clock(clock), .in1(R2872));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3078 (.out1(R3079), .clock(clock), .in1(R3078));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3280 (.out1(R3281), .clock(clock), .in1(R3280));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3527 (.out1(R3528), .clock(clock), .in1(R3527));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3719 (.out1(R3720), .clock(clock), .in1(R3719));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3907 (.out1(R3908), .clock(clock), .in1(R3907));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4140 (.out1(R4141), .clock(clock), .in1(R4140));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4318 (.out1(R4319), .clock(clock), .in1(R4318));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4492 (.out1(R4493), .clock(clock), .in1(R4492));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4711 (.out1(R4712), .clock(clock), .in1(R4711));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4875 (.out1(R4876), .clock(clock), .in1(R4875));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5035 (.out1(R5036), .clock(clock), .in1(R5035));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5240 (.out1(R5241), .clock(clock), .in1(R5240));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5390 (.out1(R5391), .clock(clock), .in1(R5390));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5536 (.out1(R5537), .clock(clock), .in1(R5536));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5727 (.out1(R5728), .clock(clock), .in1(R5727));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5863 (.out1(R5864), .clock(clock), .in1(R5863));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5995 (.out1(R5996), .clock(clock), .in1(R5995));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6171 (.out1(R6172), .clock(clock), .in1(R6171));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6292 (.out1(R6293), .clock(clock), .in1(R6292));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6409 (.out1(R6410), .clock(clock), .in1(R6409));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6572 (.out1(R6573), .clock(clock), .in1(R6572));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6679 (.out1(R6680), .clock(clock), .in1(R6679));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6782 (.out1(R6783), .clock(clock), .in1(R6782));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6930 (.out1(R6931), .clock(clock), .in1(R6930));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7023 (.out1(R7024), .clock(clock), .in1(R7023));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7112 (.out1(R7113), .clock(clock), .in1(R7112));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7246 (.out1(R7247), .clock(clock), .in1(R7246));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7325 (.out1(R7326), .clock(clock), .in1(R7325));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7400 (.out1(R7401), .clock(clock), .in1(R7400));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7520 (.out1(R7521), .clock(clock), .in1(R7520));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7585 (.out1(R7586), .clock(clock), .in1(R7585));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7646 (.out1(R7647), .clock(clock), .in1(R7646));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7752 (.out1(R7753), .clock(clock), .in1(R7752));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7803 (.out1(R7804), .clock(clock), .in1(R7803));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7850 (.out1(R7851), .clock(clock), .in1(R7850));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7942 (.out1(R7943), .clock(clock), .in1(R7942));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7979 (.out1(R7980), .clock(clock), .in1(R7979));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8012 (.out1(R8013), .clock(clock), .in1(R8012));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8090 (.out1(R8091), .clock(clock), .in1(R8090));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8113 (.out1(R8114), .clock(clock), .in1(R8113));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8132 (.out1(R8133), .clock(clock), .in1(R8132));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8195 (.out1(R8196), .clock(clock), .in1(R8195));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8240 (.out1(R8241), .clock(clock), .in1(R8240));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8259 (.out1(R8260), .clock(clock), .in1(R8259));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8270 (.out1(R8271), .clock(clock), .in1(R8270));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8281 (.out1(R8282), .clock(clock), .in1(R8281));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8292 (.out1(R8293), .clock(clock), .in1(R8292));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8303 (.out1(R8304), .clock(clock), .in1(R8303));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8314 (.out1(R8315), .clock(clock), .in1(R8314));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8325 (.out1(R8326), .clock(clock), .in1(R8325));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8336 (.out1(R8337), .clock(clock), .in1(R8336));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8347 (.out1(R8348), .clock(clock), .in1(R8347));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8372 (.out1(R8373), .clock(clock), .in1(ifout2555));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8383 (.out1(R8384), .clock(clock), .in1(ifout2466));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8394 (.out1(R8395), .clock(clock), .in1(ifout2377));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8405 (.out1(R8406), .clock(clock), .in1(ifout2288));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8416 (.out1(R8417), .clock(clock), .in1(ifout2199));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8427 (.out1(R8428), .clock(clock), .in1(ifout2110));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8438 (.out1(R8439), .clock(clock), .in1(_2502));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8439 (.out1(R8440), .clock(clock), .in1(_2416));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8440 (.out1(R8441), .clock(clock), .in1(_2330));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8441 (.out1(R8442), .clock(clock), .in1(_2244));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8442 (.out1(R8443), .clock(clock), .in1(_2158));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8443 (.out1(R8444), .clock(clock), .in1(_2072));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8444 (.out1(R8445), .clock(clock), .in1(_1980));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8445 (.out1(R8446), .clock(clock), .in1(_1970));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8446 (.out1(R8447), .clock(clock), .in1(_1964));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8447 (.out1(R8448), .clock(clock), .in1(_1952));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8448 (.out1(R8449), .clock(clock), .in1(_1946));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8449 (.out1(R8450), .clock(clock), .in1(_1936));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8450 (.out1(R8451), .clock(clock), .in1(_1894));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8451 (.out1(R8452), .clock(clock), .in1(_1884));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8452 (.out1(R8453), .clock(clock), .in1(_1878));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8453 (.out1(R8454), .clock(clock), .in1(_1866));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8454 (.out1(R8455), .clock(clock), .in1(_1860));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8455 (.out1(R8456), .clock(clock), .in1(_1850));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8456 (.out1(R8457), .clock(clock), .in1(_1808));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8457 (.out1(R8458), .clock(clock), .in1(_1798));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8458 (.out1(R8459), .clock(clock), .in1(_1792));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8459 (.out1(R8460), .clock(clock), .in1(_1780));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8460 (.out1(R8461), .clock(clock), .in1(_1774));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8461 (.out1(R8462), .clock(clock), .in1(_1764));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8462 (.out1(R8463), .clock(clock), .in1(_1722));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8463 (.out1(R8464), .clock(clock), .in1(_1712));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8464 (.out1(R8465), .clock(clock), .in1(_1706));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8465 (.out1(R8466), .clock(clock), .in1(_1694));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8466 (.out1(R8467), .clock(clock), .in1(_1688));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8467 (.out1(R8468), .clock(clock), .in1(_1678));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8468 (.out1(R8469), .clock(clock), .in1(_1636));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8469 (.out1(R8470), .clock(clock), .in1(_1626));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8470 (.out1(R8471), .clock(clock), .in1(_1620));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8471 (.out1(R8472), .clock(clock), .in1(_1608));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8472 (.out1(R8473), .clock(clock), .in1(_1602));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8473 (.out1(R8474), .clock(clock), .in1(_1592));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8474 (.out1(R8475), .clock(clock), .in1(_1550));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8475 (.out1(R8476), .clock(clock), .in1(_1540));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8476 (.out1(R8477), .clock(clock), .in1(_1534));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8477 (.out1(R8478), .clock(clock), .in1(_1522));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8478 (.out1(R8479), .clock(clock), .in1(_1516));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8479 (.out1(R8480), .clock(clock), .in1(_1506));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8480 (.out1(R8481), .clock(clock), .in1(_1464));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8481 (.out1(R8482), .clock(clock), .in1(_1454));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8482 (.out1(R8483), .clock(clock), .in1(_1448));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8483 (.out1(R8484), .clock(clock), .in1(_1436));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8484 (.out1(R8485), .clock(clock), .in1(_1430));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8485 (.out1(R8486), .clock(clock), .in1(_1420));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8486 (.out1(R8487), .clock(clock), .in1(_1378));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8487 (.out1(R8488), .clock(clock), .in1(_1368));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8488 (.out1(R8489), .clock(clock), .in1(_1362));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8489 (.out1(R8490), .clock(clock), .in1(_1350));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8490 (.out1(R8491), .clock(clock), .in1(_1344));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8491 (.out1(R8492), .clock(clock), .in1(_1334));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8492 (.out1(R8493), .clock(clock), .in1(_1292));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8493 (.out1(R8494), .clock(clock), .in1(_1282));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8494 (.out1(R8495), .clock(clock), .in1(_1276));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8495 (.out1(R8496), .clock(clock), .in1(_1264));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8496 (.out1(R8497), .clock(clock), .in1(_1258));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8497 (.out1(R8498), .clock(clock), .in1(_1248));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8498 (.out1(R8499), .clock(clock), .in1(_1987));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8499 (.out1(R8500), .clock(clock), .in1(_1901));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8500 (.out1(R8501), .clock(clock), .in1(_1815));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8501 (.out1(R8502), .clock(clock), .in1(_1729));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8502 (.out1(R8503), .clock(clock), .in1(_1643));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8503 (.out1(R8504), .clock(clock), .in1(_1557));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8504 (.out1(R8505), .clock(clock), .in1(_1471));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8505 (.out1(R8506), .clock(clock), .in1(_1385));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8506 (.out1(R8507), .clock(clock), .in1(_1299));
  SRAM op2085 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1988),.ADR(R8499));
  SRAM op1996 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1902),.ADR(R8500));
  SRAM op1907 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1816),.ADR(R8501));
  SRAM op1818 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1730),.ADR(R8502));
  SRAM op1729 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1644),.ADR(R8503));
  SRAM op1640 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1558),.ADR(R8504));
  SRAM op1551 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1472),.ADR(R8505));
  SRAM op1462 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1386),.ADR(R8506));
  SRAM op1373 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1300),.ADR(R8507));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2610 (.out1(_2495), .in1(R2873));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2600 (.out1(_2485), .in1(R2873));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2594 (.out1(_2479), .in1(R2873));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2582 (.out1(_2467), .in1(R2873));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2576 (.out1(_2461), .in1(R2873));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2566 (.out1(_2451), .in1(R2873));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2521 (.out1(_2409), .in1(R3528));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2511 (.out1(_2399), .in1(R3528));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2505 (.out1(_2393), .in1(R3528));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2493 (.out1(_2381), .in1(R3528));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2487 (.out1(_2375), .in1(R3528));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2477 (.out1(_2365), .in1(R3528));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2432 (.out1(_2323), .in1(R4141));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2422 (.out1(_2313), .in1(R4141));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2416 (.out1(_2307), .in1(R4141));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2404 (.out1(_2295), .in1(R4141));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2398 (.out1(_2289), .in1(R4141));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2388 (.out1(_2279), .in1(R4141));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2343 (.out1(_2237), .in1(R4712));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2333 (.out1(_2227), .in1(R4712));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2327 (.out1(_2221), .in1(R4712));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2315 (.out1(_2209), .in1(R4712));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2309 (.out1(_2203), .in1(R4712));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2299 (.out1(_2193), .in1(R4712));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2254 (.out1(_2151), .in1(R5241));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2244 (.out1(_2141), .in1(R5241));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2238 (.out1(_2135), .in1(R5241));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2226 (.out1(_2123), .in1(R5241));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2220 (.out1(_2117), .in1(R5241));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2210 (.out1(_2107), .in1(R5241));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2165 (.out1(_2065), .in1(R5728));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2155 (.out1(_2055), .in1(R5728));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2149 (.out1(_2049), .in1(R5728));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2137 (.out1(_2037), .in1(R5728));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2131 (.out1(_2031), .in1(R5728));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2121 (.out1(_2021), .in1(R5728));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2026 (.out1(_1929), .in1(R6172));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1937 (.out1(_1843), .in1(R6573));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1848 (.out1(_1757), .in1(R6931));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1759 (.out1(_1671), .in1(R7247));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1670 (.out1(_1585), .in1(R7521));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1581 (.out1(_1499), .in1(R7753));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1492 (.out1(_1413), .in1(R7943));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1403 (.out1(_1327), .in1(R8091));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1314 (.out1(_1241), .in1(R8196));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2611 (.out1(_2496), .in1(_2495), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2601 (.out1(_2486), .in1(_2485), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2595 (.out1(_2480), .in1(_2479), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2583 (.out1(_2468), .in1(_2467), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2577 (.out1(_2462), .in1(_2461), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2567 (.out1(_2452), .in1(_2451), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2522 (.out1(_2410), .in1(_2409), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2512 (.out1(_2400), .in1(_2399), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2506 (.out1(_2394), .in1(_2393), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2494 (.out1(_2382), .in1(_2381), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2488 (.out1(_2376), .in1(_2375), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2478 (.out1(_2366), .in1(_2365), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2433 (.out1(_2324), .in1(_2323), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2423 (.out1(_2314), .in1(_2313), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2417 (.out1(_2308), .in1(_2307), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2405 (.out1(_2296), .in1(_2295), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2399 (.out1(_2290), .in1(_2289), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2389 (.out1(_2280), .in1(_2279), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2344 (.out1(_2238), .in1(_2237), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2334 (.out1(_2228), .in1(_2227), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2328 (.out1(_2222), .in1(_2221), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2316 (.out1(_2210), .in1(_2209), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2310 (.out1(_2204), .in1(_2203), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2300 (.out1(_2194), .in1(_2193), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2255 (.out1(_2152), .in1(_2151), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2245 (.out1(_2142), .in1(_2141), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2239 (.out1(_2136), .in1(_2135), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2227 (.out1(_2124), .in1(_2123), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2221 (.out1(_2118), .in1(_2117), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2211 (.out1(_2108), .in1(_2107), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2166 (.out1(_2066), .in1(_2065), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2156 (.out1(_2056), .in1(_2055), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2150 (.out1(_2050), .in1(_2049), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2138 (.out1(_2038), .in1(_2037), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2132 (.out1(_2032), .in1(_2031), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2122 (.out1(_2022), .in1(_2021), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2027 (.out1(_1930), .in1(_1929), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1938 (.out1(_1844), .in1(_1843), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1849 (.out1(_1758), .in1(_1757), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1760 (.out1(_1672), .in1(_1671), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1671 (.out1(_1586), .in1(_1585), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1582 (.out1(_1500), .in1(_1499), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1493 (.out1(_1414), .in1(_1413), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1404 (.out1(_1328), .in1(_1327), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1315 (.out1(_1242), .in1(_1241), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2618 (.out1(_2503), .in1(b16_bitmap_2528_D), .in2(R8439));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2529 (.out1(_2417), .in1(b24_bitmap_2539_D), .in2(R8440));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2440 (.out1(_2331), .in1(b32_bitmap_2549_D), .in2(R8441));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2351 (.out1(_2245), .in1(b40_bitmap_2559_D), .in2(R8442));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2262 (.out1(_2159), .in1(b48_bitmap_2569_D), .in2(R8443));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2173 (.out1(_2073), .in1(b56_bitmap_2579_D), .in2(R8444));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2078 (.out1(_1981), .in1(b64_bitmap_2589_D), .in2(R8445));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2068 (.out1(_1971), .in1(b64_bitmap_2589_D), .in2(R8446));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2062 (.out1(_1965), .in1(b64_bitmap_2589_D), .in2(R8447));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2050 (.out1(_1953), .in1(b64_bitmap_2589_D), .in2(R8448));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2044 (.out1(_1947), .in1(b64_bitmap_2589_D), .in2(R8449));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2034 (.out1(_1937), .in1(b64_bitmap_2589_D), .in2(R8450));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1989 (.out1(_1895), .in1(b72_bitmap_2600_D), .in2(R8451));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1979 (.out1(_1885), .in1(b72_bitmap_2600_D), .in2(R8452));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1973 (.out1(_1879), .in1(b72_bitmap_2600_D), .in2(R8453));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1961 (.out1(_1867), .in1(b72_bitmap_2600_D), .in2(R8454));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1955 (.out1(_1861), .in1(b72_bitmap_2600_D), .in2(R8455));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1945 (.out1(_1851), .in1(b72_bitmap_2600_D), .in2(R8456));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1900 (.out1(_1809), .in1(b80_bitmap_2610_D), .in2(R8457));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1890 (.out1(_1799), .in1(b80_bitmap_2610_D), .in2(R8458));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1884 (.out1(_1793), .in1(b80_bitmap_2610_D), .in2(R8459));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1872 (.out1(_1781), .in1(b80_bitmap_2610_D), .in2(R8460));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1866 (.out1(_1775), .in1(b80_bitmap_2610_D), .in2(R8461));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1856 (.out1(_1765), .in1(b80_bitmap_2610_D), .in2(R8462));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1811 (.out1(_1723), .in1(b88_bitmap_2620_D), .in2(R8463));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1801 (.out1(_1713), .in1(b88_bitmap_2620_D), .in2(R8464));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1795 (.out1(_1707), .in1(b88_bitmap_2620_D), .in2(R8465));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1783 (.out1(_1695), .in1(b88_bitmap_2620_D), .in2(R8466));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1777 (.out1(_1689), .in1(b88_bitmap_2620_D), .in2(R8467));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1767 (.out1(_1679), .in1(b88_bitmap_2620_D), .in2(R8468));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1722 (.out1(_1637), .in1(b96_bitmap_2630_D), .in2(R8469));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1712 (.out1(_1627), .in1(b96_bitmap_2630_D), .in2(R8470));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1706 (.out1(_1621), .in1(b96_bitmap_2630_D), .in2(R8471));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1694 (.out1(_1609), .in1(b96_bitmap_2630_D), .in2(R8472));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1688 (.out1(_1603), .in1(b96_bitmap_2630_D), .in2(R8473));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1678 (.out1(_1593), .in1(b96_bitmap_2630_D), .in2(R8474));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1633 (.out1(_1551), .in1(b104_bitmap_2640_D), .in2(R8475));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1623 (.out1(_1541), .in1(b104_bitmap_2640_D), .in2(R8476));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1617 (.out1(_1535), .in1(b104_bitmap_2640_D), .in2(R8477));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1605 (.out1(_1523), .in1(b104_bitmap_2640_D), .in2(R8478));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1599 (.out1(_1517), .in1(b104_bitmap_2640_D), .in2(R8479));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1589 (.out1(_1507), .in1(b104_bitmap_2640_D), .in2(R8480));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1544 (.out1(_1465), .in1(b112_bitmap_2650_D), .in2(R8481));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1534 (.out1(_1455), .in1(b112_bitmap_2650_D), .in2(R8482));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1528 (.out1(_1449), .in1(b112_bitmap_2650_D), .in2(R8483));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1516 (.out1(_1437), .in1(b112_bitmap_2650_D), .in2(R8484));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1510 (.out1(_1431), .in1(b112_bitmap_2650_D), .in2(R8485));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1500 (.out1(_1421), .in1(b112_bitmap_2650_D), .in2(R8486));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1455 (.out1(_1379), .in1(b120_bitmap_2660_D), .in2(R8487));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1445 (.out1(_1369), .in1(b120_bitmap_2660_D), .in2(R8488));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1439 (.out1(_1363), .in1(b120_bitmap_2660_D), .in2(R8489));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1427 (.out1(_1351), .in1(b120_bitmap_2660_D), .in2(R8490));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1421 (.out1(_1345), .in1(b120_bitmap_2660_D), .in2(R8491));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1411 (.out1(_1335), .in1(b120_bitmap_2660_D), .in2(R8492));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1366 (.out1(_1293), .in1(b128_bitmap_2669_D), .in2(R8493));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1356 (.out1(_1283), .in1(b128_bitmap_2669_D), .in2(R8494));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1350 (.out1(_1277), .in1(b128_bitmap_2669_D), .in2(R8495));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1338 (.out1(_1265), .in1(b128_bitmap_2669_D), .in2(R8496));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1332 (.out1(_1259), .in1(b128_bitmap_2669_D), .in2(R8497));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1322 (.out1(_1249), .in1(b128_bitmap_2669_D), .in2(R8498));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2873 (.out1(R2874), .clock(clock), .in1(R2873));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3079 (.out1(R3080), .clock(clock), .in1(R3079));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3281 (.out1(R3282), .clock(clock), .in1(R3281));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3528 (.out1(R3529), .clock(clock), .in1(R3528));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3720 (.out1(R3721), .clock(clock), .in1(R3720));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3908 (.out1(R3909), .clock(clock), .in1(R3908));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4141 (.out1(R4142), .clock(clock), .in1(R4141));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4319 (.out1(R4320), .clock(clock), .in1(R4319));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4493 (.out1(R4494), .clock(clock), .in1(R4493));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4712 (.out1(R4713), .clock(clock), .in1(R4712));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4876 (.out1(R4877), .clock(clock), .in1(R4876));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5036 (.out1(R5037), .clock(clock), .in1(R5036));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5241 (.out1(R5242), .clock(clock), .in1(R5241));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5391 (.out1(R5392), .clock(clock), .in1(R5391));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5537 (.out1(R5538), .clock(clock), .in1(R5537));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5728 (.out1(R5729), .clock(clock), .in1(R5728));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5864 (.out1(R5865), .clock(clock), .in1(R5864));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5996 (.out1(R5997), .clock(clock), .in1(R5996));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6172 (.out1(R6173), .clock(clock), .in1(R6172));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6293 (.out1(R6294), .clock(clock), .in1(R6293));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6410 (.out1(R6411), .clock(clock), .in1(R6410));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6573 (.out1(R6574), .clock(clock), .in1(R6573));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6680 (.out1(R6681), .clock(clock), .in1(R6680));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6783 (.out1(R6784), .clock(clock), .in1(R6783));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6931 (.out1(R6932), .clock(clock), .in1(R6931));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7024 (.out1(R7025), .clock(clock), .in1(R7024));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7113 (.out1(R7114), .clock(clock), .in1(R7113));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7247 (.out1(R7248), .clock(clock), .in1(R7247));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7326 (.out1(R7327), .clock(clock), .in1(R7326));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7401 (.out1(R7402), .clock(clock), .in1(R7401));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7521 (.out1(R7522), .clock(clock), .in1(R7521));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7586 (.out1(R7587), .clock(clock), .in1(R7586));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7647 (.out1(R7648), .clock(clock), .in1(R7647));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7753 (.out1(R7754), .clock(clock), .in1(R7753));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7804 (.out1(R7805), .clock(clock), .in1(R7804));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7851 (.out1(R7852), .clock(clock), .in1(R7851));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7943 (.out1(R7944), .clock(clock), .in1(R7943));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7980 (.out1(R7981), .clock(clock), .in1(R7980));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8013 (.out1(R8014), .clock(clock), .in1(R8013));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8091 (.out1(R8092), .clock(clock), .in1(R8091));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8114 (.out1(R8115), .clock(clock), .in1(R8114));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8133 (.out1(R8134), .clock(clock), .in1(R8133));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8196 (.out1(R8197), .clock(clock), .in1(R8196));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8241 (.out1(R8242), .clock(clock), .in1(R8241));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8260 (.out1(R8261), .clock(clock), .in1(R8260));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8271 (.out1(R8272), .clock(clock), .in1(R8271));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8282 (.out1(R8283), .clock(clock), .in1(R8282));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8293 (.out1(R8294), .clock(clock), .in1(R8293));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8304 (.out1(R8305), .clock(clock), .in1(R8304));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8315 (.out1(R8316), .clock(clock), .in1(R8315));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8326 (.out1(R8327), .clock(clock), .in1(R8326));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8337 (.out1(R8338), .clock(clock), .in1(R8337));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8348 (.out1(R8349), .clock(clock), .in1(R8348));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8373 (.out1(R8374), .clock(clock), .in1(R8373));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8384 (.out1(R8385), .clock(clock), .in1(R8384));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8395 (.out1(R8396), .clock(clock), .in1(R8395));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8406 (.out1(R8407), .clock(clock), .in1(R8406));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8417 (.out1(R8418), .clock(clock), .in1(R8417));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8428 (.out1(R8429), .clock(clock), .in1(R8428));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8507 (.out1(R8508), .clock(clock), .in1(_1988));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8508 (.out1(R8509), .clock(clock), .in1(_1902));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8509 (.out1(R8510), .clock(clock), .in1(_1816));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8510 (.out1(R8511), .clock(clock), .in1(_1730));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8511 (.out1(R8512), .clock(clock), .in1(_1644));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8512 (.out1(R8513), .clock(clock), .in1(_1558));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8513 (.out1(R8514), .clock(clock), .in1(_1472));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8514 (.out1(R8515), .clock(clock), .in1(_1386));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8515 (.out1(R8516), .clock(clock), .in1(_1300));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8516 (.out1(R8517), .clock(clock), .in1(_2496));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8517 (.out1(R8518), .clock(clock), .in1(_2486));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8518 (.out1(R8519), .clock(clock), .in1(_2480));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8519 (.out1(R8520), .clock(clock), .in1(_2468));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8520 (.out1(R8521), .clock(clock), .in1(_2462));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8521 (.out1(R8522), .clock(clock), .in1(_2452));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8522 (.out1(R8523), .clock(clock), .in1(_2410));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8523 (.out1(R8524), .clock(clock), .in1(_2400));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8524 (.out1(R8525), .clock(clock), .in1(_2394));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8525 (.out1(R8526), .clock(clock), .in1(_2382));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8526 (.out1(R8527), .clock(clock), .in1(_2376));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8527 (.out1(R8528), .clock(clock), .in1(_2366));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8528 (.out1(R8529), .clock(clock), .in1(_2324));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8529 (.out1(R8530), .clock(clock), .in1(_2314));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8530 (.out1(R8531), .clock(clock), .in1(_2308));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8531 (.out1(R8532), .clock(clock), .in1(_2296));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8532 (.out1(R8533), .clock(clock), .in1(_2290));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8533 (.out1(R8534), .clock(clock), .in1(_2280));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8534 (.out1(R8535), .clock(clock), .in1(_2238));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8535 (.out1(R8536), .clock(clock), .in1(_2228));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8536 (.out1(R8537), .clock(clock), .in1(_2222));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8537 (.out1(R8538), .clock(clock), .in1(_2210));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8538 (.out1(R8539), .clock(clock), .in1(_2204));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8539 (.out1(R8540), .clock(clock), .in1(_2194));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8540 (.out1(R8541), .clock(clock), .in1(_2152));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8541 (.out1(R8542), .clock(clock), .in1(_2142));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8542 (.out1(R8543), .clock(clock), .in1(_2136));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8543 (.out1(R8544), .clock(clock), .in1(_2124));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8544 (.out1(R8545), .clock(clock), .in1(_2118));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8545 (.out1(R8546), .clock(clock), .in1(_2108));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8546 (.out1(R8547), .clock(clock), .in1(_2066));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8547 (.out1(R8548), .clock(clock), .in1(_2056));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8548 (.out1(R8549), .clock(clock), .in1(_2050));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8549 (.out1(R8550), .clock(clock), .in1(_2038));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8550 (.out1(R8551), .clock(clock), .in1(_2032));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8551 (.out1(R8552), .clock(clock), .in1(_2022));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8552 (.out1(R8553), .clock(clock), .in1(_1930));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8553 (.out1(R8554), .clock(clock), .in1(_1844));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8554 (.out1(R8555), .clock(clock), .in1(_1758));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8555 (.out1(R8556), .clock(clock), .in1(_1672));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8556 (.out1(R8557), .clock(clock), .in1(_1586));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8557 (.out1(R8558), .clock(clock), .in1(_1500));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8558 (.out1(R8559), .clock(clock), .in1(_1414));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8559 (.out1(R8560), .clock(clock), .in1(_1328));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8560 (.out1(R8561), .clock(clock), .in1(_1242));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8561 (.out1(R8562), .clock(clock), .in1(_2503));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8562 (.out1(R8563), .clock(clock), .in1(_2417));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8563 (.out1(R8564), .clock(clock), .in1(_2331));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8564 (.out1(R8565), .clock(clock), .in1(_2245));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8565 (.out1(R8566), .clock(clock), .in1(_2159));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8566 (.out1(R8567), .clock(clock), .in1(_2073));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8567 (.out1(R8568), .clock(clock), .in1(_1981));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8568 (.out1(R8569), .clock(clock), .in1(_1971));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8569 (.out1(R8570), .clock(clock), .in1(_1965));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8570 (.out1(R8571), .clock(clock), .in1(_1953));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8571 (.out1(R8572), .clock(clock), .in1(_1947));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8572 (.out1(R8573), .clock(clock), .in1(_1937));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8573 (.out1(R8574), .clock(clock), .in1(_1895));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8574 (.out1(R8575), .clock(clock), .in1(_1885));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8575 (.out1(R8576), .clock(clock), .in1(_1879));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8576 (.out1(R8577), .clock(clock), .in1(_1867));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8577 (.out1(R8578), .clock(clock), .in1(_1861));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8578 (.out1(R8579), .clock(clock), .in1(_1851));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8579 (.out1(R8580), .clock(clock), .in1(_1809));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8580 (.out1(R8581), .clock(clock), .in1(_1799));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8581 (.out1(R8582), .clock(clock), .in1(_1793));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8582 (.out1(R8583), .clock(clock), .in1(_1781));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8583 (.out1(R8584), .clock(clock), .in1(_1775));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8584 (.out1(R8585), .clock(clock), .in1(_1765));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8585 (.out1(R8586), .clock(clock), .in1(_1723));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8586 (.out1(R8587), .clock(clock), .in1(_1713));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8587 (.out1(R8588), .clock(clock), .in1(_1707));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8588 (.out1(R8589), .clock(clock), .in1(_1695));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8589 (.out1(R8590), .clock(clock), .in1(_1689));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8590 (.out1(R8591), .clock(clock), .in1(_1679));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8591 (.out1(R8592), .clock(clock), .in1(_1637));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8592 (.out1(R8593), .clock(clock), .in1(_1627));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8593 (.out1(R8594), .clock(clock), .in1(_1621));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8594 (.out1(R8595), .clock(clock), .in1(_1609));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8595 (.out1(R8596), .clock(clock), .in1(_1603));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8596 (.out1(R8597), .clock(clock), .in1(_1593));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8597 (.out1(R8598), .clock(clock), .in1(_1551));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8598 (.out1(R8599), .clock(clock), .in1(_1541));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8599 (.out1(R8600), .clock(clock), .in1(_1535));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8600 (.out1(R8601), .clock(clock), .in1(_1523));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8601 (.out1(R8602), .clock(clock), .in1(_1517));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8602 (.out1(R8603), .clock(clock), .in1(_1507));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8603 (.out1(R8604), .clock(clock), .in1(_1465));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8604 (.out1(R8605), .clock(clock), .in1(_1455));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8605 (.out1(R8606), .clock(clock), .in1(_1449));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8606 (.out1(R8607), .clock(clock), .in1(_1437));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8607 (.out1(R8608), .clock(clock), .in1(_1431));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8608 (.out1(R8609), .clock(clock), .in1(_1421));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8609 (.out1(R8610), .clock(clock), .in1(_1379));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8610 (.out1(R8611), .clock(clock), .in1(_1369));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8611 (.out1(R8612), .clock(clock), .in1(_1363));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8612 (.out1(R8613), .clock(clock), .in1(_1351));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8613 (.out1(R8614), .clock(clock), .in1(_1345));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8614 (.out1(R8615), .clock(clock), .in1(_1335));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8615 (.out1(R8616), .clock(clock), .in1(_1293));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8616 (.out1(R8617), .clock(clock), .in1(_1283));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8617 (.out1(R8618), .clock(clock), .in1(_1277));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8618 (.out1(R8619), .clock(clock), .in1(_1265));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8619 (.out1(R8620), .clock(clock), .in1(_1259));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8620 (.out1(R8621), .clock(clock), .in1(_1249));
  SRAM op2619 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2504),.ADR(R8562));
  SRAM op2530 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2418),.ADR(R8563));
  SRAM op2441 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2332),.ADR(R8564));
  SRAM op2352 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2246),.ADR(R8565));
  SRAM op2263 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2160),.ADR(R8566));
  SRAM op2174 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2074),.ADR(R8567));
  SRAM op2079 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1982),.ADR(R8568));
  SRAM op2069 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1972),.ADR(R8569));
  SRAM op2063 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1966),.ADR(R8570));
  SRAM op2051 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1954),.ADR(R8571));
  SRAM op2045 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1948),.ADR(R8572));
  SRAM op2035 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1938),.ADR(R8573));
  SRAM op1990 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1896),.ADR(R8574));
  SRAM op1980 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1886),.ADR(R8575));
  SRAM op1974 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1880),.ADR(R8576));
  SRAM op1962 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1868),.ADR(R8577));
  SRAM op1956 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1862),.ADR(R8578));
  SRAM op1946 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1852),.ADR(R8579));
  SRAM op1901 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1810),.ADR(R8580));
  SRAM op1891 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1800),.ADR(R8581));
  SRAM op1885 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1794),.ADR(R8582));
  SRAM op1873 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1782),.ADR(R8583));
  SRAM op1867 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1776),.ADR(R8584));
  SRAM op1857 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1766),.ADR(R8585));
  SRAM op1812 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1724),.ADR(R8586));
  SRAM op1802 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1714),.ADR(R8587));
  SRAM op1796 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1708),.ADR(R8588));
  SRAM op1784 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1696),.ADR(R8589));
  SRAM op1778 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1690),.ADR(R8590));
  SRAM op1768 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1680),.ADR(R8591));
  SRAM op1723 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1638),.ADR(R8592));
  SRAM op1713 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1628),.ADR(R8593));
  SRAM op1707 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1622),.ADR(R8594));
  SRAM op1695 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1610),.ADR(R8595));
  SRAM op1689 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1604),.ADR(R8596));
  SRAM op1679 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1594),.ADR(R8597));
  SRAM op1634 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1552),.ADR(R8598));
  SRAM op1624 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1542),.ADR(R8599));
  SRAM op1618 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1536),.ADR(R8600));
  SRAM op1606 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1524),.ADR(R8601));
  SRAM op1600 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1518),.ADR(R8602));
  SRAM op1590 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1508),.ADR(R8603));
  SRAM op1545 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1466),.ADR(R8604));
  SRAM op1535 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1456),.ADR(R8605));
  SRAM op1529 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1450),.ADR(R8606));
  SRAM op1517 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1438),.ADR(R8607));
  SRAM op1511 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1432),.ADR(R8608));
  SRAM op1501 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1422),.ADR(R8609));
  SRAM op1456 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1380),.ADR(R8610));
  SRAM op1446 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1370),.ADR(R8611));
  SRAM op1440 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1364),.ADR(R8612));
  SRAM op1428 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1352),.ADR(R8613));
  SRAM op1422 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1346),.ADR(R8614));
  SRAM op1412 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1336),.ADR(R8615));
  SRAM op1367 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1294),.ADR(R8616));
  SRAM op1357 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1284),.ADR(R8617));
  SRAM op1351 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1278),.ADR(R8618));
  SRAM op1339 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1266),.ADR(R8619));
  SRAM op1333 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1260),.ADR(R8620));
  SRAM op1323 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1250),.ADR(R8621));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2560 (.out1(_2445), .in1(R2874));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2471 (.out1(_2359), .in1(R3529));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2382 (.out1(_2273), .in1(R4142));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2293 (.out1(_2187), .in1(R4713));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2204 (.out1(_2101), .in1(R5242));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2115 (.out1(_2015), .in1(R5729));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2086 (.out1(_1989), .in1(7 'd 64), .in2(R6294));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1997 (.out1(_1903), .in1(7 'd 64), .in2(R6681));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1908 (.out1(_1817), .in1(7 'd 64), .in2(R7025));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1819 (.out1(_1731), .in1(7 'd 64), .in2(R7327));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1730 (.out1(_1645), .in1(7 'd 64), .in2(R7587));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1641 (.out1(_1559), .in1(7 'd 64), .in2(R7805));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1552 (.out1(_1473), .in1(7 'd 64), .in2(R7981));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1463 (.out1(_1387), .in1(7 'd 64), .in2(R8115));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1374 (.out1(_1301), .in1(7 'd 64), .in2(R8242));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2561 (.out1(_2446), .in1(_2445), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2472 (.out1(_2360), .in1(_2359), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2383 (.out1(_2274), .in1(_2273), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2294 (.out1(_2188), .in1(_2187), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2205 (.out1(_2102), .in1(_2101), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2116 (.out1(_2016), .in1(_2015), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2612 (.out1(_2497), .in1(b16_bitmap_2528_D), .in2(R8517));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2602 (.out1(_2487), .in1(b16_bitmap_2528_D), .in2(R8518));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2596 (.out1(_2481), .in1(b16_bitmap_2528_D), .in2(R8519));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2584 (.out1(_2469), .in1(b16_bitmap_2528_D), .in2(R8520));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2578 (.out1(_2463), .in1(b16_bitmap_2528_D), .in2(R8521));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2568 (.out1(_2453), .in1(b16_bitmap_2528_D), .in2(R8522));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2523 (.out1(_2411), .in1(b24_bitmap_2539_D), .in2(R8523));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2513 (.out1(_2401), .in1(b24_bitmap_2539_D), .in2(R8524));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2507 (.out1(_2395), .in1(b24_bitmap_2539_D), .in2(R8525));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2495 (.out1(_2383), .in1(b24_bitmap_2539_D), .in2(R8526));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2489 (.out1(_2377), .in1(b24_bitmap_2539_D), .in2(R8527));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2479 (.out1(_2367), .in1(b24_bitmap_2539_D), .in2(R8528));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2434 (.out1(_2325), .in1(b32_bitmap_2549_D), .in2(R8529));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2424 (.out1(_2315), .in1(b32_bitmap_2549_D), .in2(R8530));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2418 (.out1(_2309), .in1(b32_bitmap_2549_D), .in2(R8531));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2406 (.out1(_2297), .in1(b32_bitmap_2549_D), .in2(R8532));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2400 (.out1(_2291), .in1(b32_bitmap_2549_D), .in2(R8533));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2390 (.out1(_2281), .in1(b32_bitmap_2549_D), .in2(R8534));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2345 (.out1(_2239), .in1(b40_bitmap_2559_D), .in2(R8535));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2335 (.out1(_2229), .in1(b40_bitmap_2559_D), .in2(R8536));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2329 (.out1(_2223), .in1(b40_bitmap_2559_D), .in2(R8537));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2317 (.out1(_2211), .in1(b40_bitmap_2559_D), .in2(R8538));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2311 (.out1(_2205), .in1(b40_bitmap_2559_D), .in2(R8539));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2301 (.out1(_2195), .in1(b40_bitmap_2559_D), .in2(R8540));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2256 (.out1(_2153), .in1(b48_bitmap_2569_D), .in2(R8541));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2246 (.out1(_2143), .in1(b48_bitmap_2569_D), .in2(R8542));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2240 (.out1(_2137), .in1(b48_bitmap_2569_D), .in2(R8543));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2228 (.out1(_2125), .in1(b48_bitmap_2569_D), .in2(R8544));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2222 (.out1(_2119), .in1(b48_bitmap_2569_D), .in2(R8545));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2212 (.out1(_2109), .in1(b48_bitmap_2569_D), .in2(R8546));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2167 (.out1(_2067), .in1(b56_bitmap_2579_D), .in2(R8547));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2157 (.out1(_2057), .in1(b56_bitmap_2579_D), .in2(R8548));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2151 (.out1(_2051), .in1(b56_bitmap_2579_D), .in2(R8549));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2139 (.out1(_2039), .in1(b56_bitmap_2579_D), .in2(R8550));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2133 (.out1(_2033), .in1(b56_bitmap_2579_D), .in2(R8551));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2123 (.out1(_2023), .in1(b56_bitmap_2579_D), .in2(R8552));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2028 (.out1(_1931), .in1(b64_bitmap_2589_D), .in2(R8553));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1939 (.out1(_1845), .in1(b72_bitmap_2600_D), .in2(R8554));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1850 (.out1(_1759), .in1(b80_bitmap_2610_D), .in2(R8555));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1761 (.out1(_1673), .in1(b88_bitmap_2620_D), .in2(R8556));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1672 (.out1(_1587), .in1(b96_bitmap_2630_D), .in2(R8557));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1583 (.out1(_1501), .in1(b104_bitmap_2640_D), .in2(R8558));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1494 (.out1(_1415), .in1(b112_bitmap_2650_D), .in2(R8559));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1405 (.out1(_1329), .in1(b120_bitmap_2660_D), .in2(R8560));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1316 (.out1(_1243), .in1(b128_bitmap_2669_D), .in2(R8561));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2087 (.out1(_1990), .in1(R8508), .in2(_1989));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2080 (.out1(_1983), .in1(7 'd 64), .in2(R6294));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2070 (.out1(_1973), .in1(7 'd 64), .in2(R6294));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2052 (.out1(_1955), .in1(7 'd 64), .in2(R6294));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1998 (.out1(_1904), .in1(R8509), .in2(_1903));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1991 (.out1(_1897), .in1(7 'd 64), .in2(R6681));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1981 (.out1(_1887), .in1(7 'd 64), .in2(R6681));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1963 (.out1(_1869), .in1(7 'd 64), .in2(R6681));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1909 (.out1(_1818), .in1(R8510), .in2(_1817));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1902 (.out1(_1811), .in1(7 'd 64), .in2(R7025));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1892 (.out1(_1801), .in1(7 'd 64), .in2(R7025));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1874 (.out1(_1783), .in1(7 'd 64), .in2(R7025));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1820 (.out1(_1732), .in1(R8511), .in2(_1731));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1813 (.out1(_1725), .in1(7 'd 64), .in2(R7327));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1803 (.out1(_1715), .in1(7 'd 64), .in2(R7327));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1785 (.out1(_1697), .in1(7 'd 64), .in2(R7327));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1731 (.out1(_1646), .in1(R8512), .in2(_1645));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1724 (.out1(_1639), .in1(7 'd 64), .in2(R7587));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1714 (.out1(_1629), .in1(7 'd 64), .in2(R7587));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1696 (.out1(_1611), .in1(7 'd 64), .in2(R7587));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1642 (.out1(_1560), .in1(R8513), .in2(_1559));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1635 (.out1(_1553), .in1(7 'd 64), .in2(R7805));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1625 (.out1(_1543), .in1(7 'd 64), .in2(R7805));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1607 (.out1(_1525), .in1(7 'd 64), .in2(R7805));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1553 (.out1(_1474), .in1(R8514), .in2(_1473));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1546 (.out1(_1467), .in1(7 'd 64), .in2(R7981));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1536 (.out1(_1457), .in1(7 'd 64), .in2(R7981));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1518 (.out1(_1439), .in1(7 'd 64), .in2(R7981));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1464 (.out1(_1388), .in1(R8515), .in2(_1387));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1457 (.out1(_1381), .in1(7 'd 64), .in2(R8115));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1447 (.out1(_1371), .in1(7 'd 64), .in2(R8115));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1429 (.out1(_1353), .in1(7 'd 64), .in2(R8115));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1375 (.out1(_1302), .in1(R8516), .in2(_1301));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1368 (.out1(_1295), .in1(7 'd 64), .in2(R8242));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1358 (.out1(_1285), .in1(7 'd 64), .in2(R8242));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1340 (.out1(_1267), .in1(7 'd 64), .in2(R8242));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2874 (.out1(R2875), .clock(clock), .in1(R2874));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3080 (.out1(R3081), .clock(clock), .in1(R3080));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3282 (.out1(R3283), .clock(clock), .in1(R3282));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3529 (.out1(R3530), .clock(clock), .in1(R3529));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3721 (.out1(R3722), .clock(clock), .in1(R3721));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3909 (.out1(R3910), .clock(clock), .in1(R3909));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4142 (.out1(R4143), .clock(clock), .in1(R4142));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4320 (.out1(R4321), .clock(clock), .in1(R4320));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4494 (.out1(R4495), .clock(clock), .in1(R4494));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4713 (.out1(R4714), .clock(clock), .in1(R4713));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4877 (.out1(R4878), .clock(clock), .in1(R4877));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5037 (.out1(R5038), .clock(clock), .in1(R5037));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5242 (.out1(R5243), .clock(clock), .in1(R5242));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5392 (.out1(R5393), .clock(clock), .in1(R5392));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5538 (.out1(R5539), .clock(clock), .in1(R5538));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5729 (.out1(R5730), .clock(clock), .in1(R5729));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5865 (.out1(R5866), .clock(clock), .in1(R5865));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5997 (.out1(R5998), .clock(clock), .in1(R5997));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6173 (.out1(R6174), .clock(clock), .in1(R6173));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6294 (.out1(R6295), .clock(clock), .in1(R6294));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6411 (.out1(R6412), .clock(clock), .in1(R6411));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6574 (.out1(R6575), .clock(clock), .in1(R6574));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6681 (.out1(R6682), .clock(clock), .in1(R6681));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6784 (.out1(R6785), .clock(clock), .in1(R6784));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6932 (.out1(R6933), .clock(clock), .in1(R6932));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7025 (.out1(R7026), .clock(clock), .in1(R7025));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7114 (.out1(R7115), .clock(clock), .in1(R7114));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7248 (.out1(R7249), .clock(clock), .in1(R7248));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7327 (.out1(R7328), .clock(clock), .in1(R7327));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7402 (.out1(R7403), .clock(clock), .in1(R7402));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7522 (.out1(R7523), .clock(clock), .in1(R7522));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7587 (.out1(R7588), .clock(clock), .in1(R7587));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7648 (.out1(R7649), .clock(clock), .in1(R7648));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7754 (.out1(R7755), .clock(clock), .in1(R7754));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7805 (.out1(R7806), .clock(clock), .in1(R7805));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7852 (.out1(R7853), .clock(clock), .in1(R7852));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7944 (.out1(R7945), .clock(clock), .in1(R7944));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7981 (.out1(R7982), .clock(clock), .in1(R7981));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8014 (.out1(R8015), .clock(clock), .in1(R8014));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8092 (.out1(R8093), .clock(clock), .in1(R8092));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8115 (.out1(R8116), .clock(clock), .in1(R8115));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8134 (.out1(R8135), .clock(clock), .in1(R8134));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8197 (.out1(R8198), .clock(clock), .in1(R8197));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8242 (.out1(R8243), .clock(clock), .in1(R8242));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8261 (.out1(R8262), .clock(clock), .in1(R8261));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8272 (.out1(R8273), .clock(clock), .in1(R8272));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8283 (.out1(R8284), .clock(clock), .in1(R8283));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8294 (.out1(R8295), .clock(clock), .in1(R8294));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8305 (.out1(R8306), .clock(clock), .in1(R8305));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8316 (.out1(R8317), .clock(clock), .in1(R8316));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8327 (.out1(R8328), .clock(clock), .in1(R8327));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8338 (.out1(R8339), .clock(clock), .in1(R8338));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8349 (.out1(R8350), .clock(clock), .in1(R8349));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8374 (.out1(R8375), .clock(clock), .in1(R8374));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8385 (.out1(R8386), .clock(clock), .in1(R8385));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8396 (.out1(R8397), .clock(clock), .in1(R8396));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8407 (.out1(R8408), .clock(clock), .in1(R8407));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8418 (.out1(R8419), .clock(clock), .in1(R8418));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8429 (.out1(R8430), .clock(clock), .in1(R8429));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8621 (.out1(R8622), .clock(clock), .in1(_2504));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8622 (.out1(R8623), .clock(clock), .in1(_2418));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8623 (.out1(R8624), .clock(clock), .in1(_2332));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8624 (.out1(R8625), .clock(clock), .in1(_2246));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8625 (.out1(R8626), .clock(clock), .in1(_2160));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8626 (.out1(R8627), .clock(clock), .in1(_2074));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8627 (.out1(R8628), .clock(clock), .in1(_1982));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8628 (.out1(R8629), .clock(clock), .in1(_1972));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8629 (.out1(R8630), .clock(clock), .in1(_1966));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8630 (.out1(R8631), .clock(clock), .in1(_1954));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8631 (.out1(R8632), .clock(clock), .in1(_1948));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8632 (.out1(R8633), .clock(clock), .in1(_1938));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8633 (.out1(R8634), .clock(clock), .in1(_1896));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8634 (.out1(R8635), .clock(clock), .in1(_1886));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8635 (.out1(R8636), .clock(clock), .in1(_1880));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8636 (.out1(R8637), .clock(clock), .in1(_1868));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8637 (.out1(R8638), .clock(clock), .in1(_1862));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8638 (.out1(R8639), .clock(clock), .in1(_1852));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8639 (.out1(R8640), .clock(clock), .in1(_1810));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8640 (.out1(R8641), .clock(clock), .in1(_1800));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8641 (.out1(R8642), .clock(clock), .in1(_1794));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8642 (.out1(R8643), .clock(clock), .in1(_1782));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8643 (.out1(R8644), .clock(clock), .in1(_1776));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8644 (.out1(R8645), .clock(clock), .in1(_1766));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8645 (.out1(R8646), .clock(clock), .in1(_1724));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8646 (.out1(R8647), .clock(clock), .in1(_1714));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8647 (.out1(R8648), .clock(clock), .in1(_1708));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8648 (.out1(R8649), .clock(clock), .in1(_1696));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8649 (.out1(R8650), .clock(clock), .in1(_1690));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8650 (.out1(R8651), .clock(clock), .in1(_1680));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8651 (.out1(R8652), .clock(clock), .in1(_1638));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8652 (.out1(R8653), .clock(clock), .in1(_1628));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8653 (.out1(R8654), .clock(clock), .in1(_1622));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8654 (.out1(R8655), .clock(clock), .in1(_1610));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8655 (.out1(R8656), .clock(clock), .in1(_1604));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8656 (.out1(R8657), .clock(clock), .in1(_1594));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8657 (.out1(R8658), .clock(clock), .in1(_1552));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8658 (.out1(R8659), .clock(clock), .in1(_1542));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8659 (.out1(R8660), .clock(clock), .in1(_1536));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8660 (.out1(R8661), .clock(clock), .in1(_1524));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8661 (.out1(R8662), .clock(clock), .in1(_1518));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8662 (.out1(R8663), .clock(clock), .in1(_1508));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8663 (.out1(R8664), .clock(clock), .in1(_1466));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8664 (.out1(R8665), .clock(clock), .in1(_1456));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8665 (.out1(R8666), .clock(clock), .in1(_1450));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8666 (.out1(R8667), .clock(clock), .in1(_1438));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8667 (.out1(R8668), .clock(clock), .in1(_1432));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8668 (.out1(R8669), .clock(clock), .in1(_1422));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8669 (.out1(R8670), .clock(clock), .in1(_1380));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8670 (.out1(R8671), .clock(clock), .in1(_1370));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8671 (.out1(R8672), .clock(clock), .in1(_1364));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8672 (.out1(R8673), .clock(clock), .in1(_1352));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8673 (.out1(R8674), .clock(clock), .in1(_1346));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8674 (.out1(R8675), .clock(clock), .in1(_1336));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8675 (.out1(R8676), .clock(clock), .in1(_1294));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8676 (.out1(R8677), .clock(clock), .in1(_1284));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8677 (.out1(R8678), .clock(clock), .in1(_1278));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8678 (.out1(R8679), .clock(clock), .in1(_1266));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8679 (.out1(R8680), .clock(clock), .in1(_1260));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8680 (.out1(R8681), .clock(clock), .in1(_1250));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8681 (.out1(R8682), .clock(clock), .in1(_2446));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8682 (.out1(R8683), .clock(clock), .in1(_2360));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8683 (.out1(R8684), .clock(clock), .in1(_2274));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8684 (.out1(R8685), .clock(clock), .in1(_2188));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8685 (.out1(R8686), .clock(clock), .in1(_2102));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8686 (.out1(R8687), .clock(clock), .in1(_2016));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8687 (.out1(R8688), .clock(clock), .in1(_2497));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8688 (.out1(R8689), .clock(clock), .in1(_2487));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8689 (.out1(R8690), .clock(clock), .in1(_2481));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8690 (.out1(R8691), .clock(clock), .in1(_2469));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8691 (.out1(R8692), .clock(clock), .in1(_2463));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8692 (.out1(R8693), .clock(clock), .in1(_2453));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8693 (.out1(R8694), .clock(clock), .in1(_2411));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8694 (.out1(R8695), .clock(clock), .in1(_2401));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8695 (.out1(R8696), .clock(clock), .in1(_2395));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8696 (.out1(R8697), .clock(clock), .in1(_2383));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8697 (.out1(R8698), .clock(clock), .in1(_2377));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8698 (.out1(R8699), .clock(clock), .in1(_2367));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8699 (.out1(R8700), .clock(clock), .in1(_2325));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8700 (.out1(R8701), .clock(clock), .in1(_2315));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8701 (.out1(R8702), .clock(clock), .in1(_2309));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8702 (.out1(R8703), .clock(clock), .in1(_2297));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8703 (.out1(R8704), .clock(clock), .in1(_2291));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8704 (.out1(R8705), .clock(clock), .in1(_2281));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8705 (.out1(R8706), .clock(clock), .in1(_2239));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8706 (.out1(R8707), .clock(clock), .in1(_2229));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8707 (.out1(R8708), .clock(clock), .in1(_2223));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8708 (.out1(R8709), .clock(clock), .in1(_2211));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8709 (.out1(R8710), .clock(clock), .in1(_2205));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8710 (.out1(R8711), .clock(clock), .in1(_2195));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8711 (.out1(R8712), .clock(clock), .in1(_2153));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8712 (.out1(R8713), .clock(clock), .in1(_2143));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8713 (.out1(R8714), .clock(clock), .in1(_2137));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8714 (.out1(R8715), .clock(clock), .in1(_2125));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8715 (.out1(R8716), .clock(clock), .in1(_2119));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8716 (.out1(R8717), .clock(clock), .in1(_2109));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8717 (.out1(R8718), .clock(clock), .in1(_2067));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8718 (.out1(R8719), .clock(clock), .in1(_2057));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8719 (.out1(R8720), .clock(clock), .in1(_2051));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8720 (.out1(R8721), .clock(clock), .in1(_2039));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8721 (.out1(R8722), .clock(clock), .in1(_2033));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8722 (.out1(R8723), .clock(clock), .in1(_2023));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8723 (.out1(R8724), .clock(clock), .in1(_1931));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8724 (.out1(R8725), .clock(clock), .in1(_1845));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8725 (.out1(R8726), .clock(clock), .in1(_1759));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8726 (.out1(R8727), .clock(clock), .in1(_1673));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8727 (.out1(R8728), .clock(clock), .in1(_1587));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8728 (.out1(R8729), .clock(clock), .in1(_1501));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8729 (.out1(R8730), .clock(clock), .in1(_1415));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8730 (.out1(R8731), .clock(clock), .in1(_1329));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8731 (.out1(R8732), .clock(clock), .in1(_1243));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8732 (.out1(R8733), .clock(clock), .in1(_1990));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8733 (.out1(R8734), .clock(clock), .in1(_1983));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8734 (.out1(R8735), .clock(clock), .in1(_1973));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8735 (.out1(R8736), .clock(clock), .in1(_1955));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8736 (.out1(R8737), .clock(clock), .in1(_1904));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8737 (.out1(R8738), .clock(clock), .in1(_1897));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8738 (.out1(R8739), .clock(clock), .in1(_1887));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8739 (.out1(R8740), .clock(clock), .in1(_1869));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8740 (.out1(R8741), .clock(clock), .in1(_1818));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8741 (.out1(R8742), .clock(clock), .in1(_1811));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8742 (.out1(R8743), .clock(clock), .in1(_1801));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8743 (.out1(R8744), .clock(clock), .in1(_1783));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8744 (.out1(R8745), .clock(clock), .in1(_1732));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8745 (.out1(R8746), .clock(clock), .in1(_1725));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8746 (.out1(R8747), .clock(clock), .in1(_1715));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8747 (.out1(R8748), .clock(clock), .in1(_1697));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8748 (.out1(R8749), .clock(clock), .in1(_1646));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8749 (.out1(R8750), .clock(clock), .in1(_1639));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8750 (.out1(R8751), .clock(clock), .in1(_1629));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8751 (.out1(R8752), .clock(clock), .in1(_1611));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8752 (.out1(R8753), .clock(clock), .in1(_1560));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8753 (.out1(R8754), .clock(clock), .in1(_1553));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8754 (.out1(R8755), .clock(clock), .in1(_1543));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8755 (.out1(R8756), .clock(clock), .in1(_1525));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8756 (.out1(R8757), .clock(clock), .in1(_1474));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8757 (.out1(R8758), .clock(clock), .in1(_1467));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8758 (.out1(R8759), .clock(clock), .in1(_1457));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8759 (.out1(R8760), .clock(clock), .in1(_1439));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8760 (.out1(R8761), .clock(clock), .in1(_1388));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8761 (.out1(R8762), .clock(clock), .in1(_1381));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8762 (.out1(R8763), .clock(clock), .in1(_1371));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8763 (.out1(R8764), .clock(clock), .in1(_1353));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8764 (.out1(R8765), .clock(clock), .in1(_1302));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8765 (.out1(R8766), .clock(clock), .in1(_1295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8766 (.out1(R8767), .clock(clock), .in1(_1285));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8767 (.out1(R8768), .clock(clock), .in1(_1267));
  SRAM op2613 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2498),.ADR(R8688));
  SRAM op2603 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2488),.ADR(R8689));
  SRAM op2597 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2482),.ADR(R8690));
  SRAM op2585 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2470),.ADR(R8691));
  SRAM op2579 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2464),.ADR(R8692));
  SRAM op2569 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2454),.ADR(R8693));
  SRAM op2524 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2412),.ADR(R8694));
  SRAM op2514 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2402),.ADR(R8695));
  SRAM op2508 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2396),.ADR(R8696));
  SRAM op2496 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2384),.ADR(R8697));
  SRAM op2490 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2378),.ADR(R8698));
  SRAM op2480 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2368),.ADR(R8699));
  SRAM op2435 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2326),.ADR(R8700));
  SRAM op2425 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2316),.ADR(R8701));
  SRAM op2419 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2310),.ADR(R8702));
  SRAM op2407 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2298),.ADR(R8703));
  SRAM op2401 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2292),.ADR(R8704));
  SRAM op2391 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2282),.ADR(R8705));
  SRAM op2346 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2240),.ADR(R8706));
  SRAM op2336 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2230),.ADR(R8707));
  SRAM op2330 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2224),.ADR(R8708));
  SRAM op2318 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2212),.ADR(R8709));
  SRAM op2312 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2206),.ADR(R8710));
  SRAM op2302 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2196),.ADR(R8711));
  SRAM op2257 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2154),.ADR(R8712));
  SRAM op2247 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2144),.ADR(R8713));
  SRAM op2241 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2138),.ADR(R8714));
  SRAM op2229 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2126),.ADR(R8715));
  SRAM op2223 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2120),.ADR(R8716));
  SRAM op2213 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2110),.ADR(R8717));
  SRAM op2168 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2068),.ADR(R8718));
  SRAM op2158 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2058),.ADR(R8719));
  SRAM op2152 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2052),.ADR(R8720));
  SRAM op2140 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2040),.ADR(R8721));
  SRAM op2134 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2034),.ADR(R8722));
  SRAM op2124 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2024),.ADR(R8723));
  SRAM op2029 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1932),.ADR(R8724));
  SRAM op1940 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1846),.ADR(R8725));
  SRAM op1851 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1760),.ADR(R8726));
  SRAM op1762 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1674),.ADR(R8727));
  SRAM op1673 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1588),.ADR(R8728));
  SRAM op1584 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1502),.ADR(R8729));
  SRAM op1495 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1416),.ADR(R8730));
  SRAM op1406 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1330),.ADR(R8731));
  SRAM op1317 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1244),.ADR(R8732));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2088 (.out1(_1991), .in1(R8733), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1999 (.out1(_1905), .in1(R8737), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1910 (.out1(_1819), .in1(R8741), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1821 (.out1(_1733), .in1(R8745), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1732 (.out1(_1647), .in1(R8749), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1643 (.out1(_1561), .in1(R8753), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1554 (.out1(_1475), .in1(R8757), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1465 (.out1(_1389), .in1(R8761), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1376 (.out1(_1303), .in1(R8765), .in2(1 'd 1));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2620 (.out1(_2505), .in1(7 'd 64), .in2(R3081));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2531 (.out1(_2419), .in1(7 'd 64), .in2(R3722));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2442 (.out1(_2333), .in1(7 'd 64), .in2(R4321));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2353 (.out1(_2247), .in1(7 'd 64), .in2(R4878));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2264 (.out1(_2161), .in1(7 'd 64), .in2(R5393));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2175 (.out1(_2075), .in1(7 'd 64), .in2(R5866));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2081 (.out1(_1984), .in1(R8628), .in2(R8734));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2071 (.out1(_1974), .in1(R8629), .in2(R8735));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2064 (.out1(_1967), .in1(7 'd 64), .in2(R6295));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2053 (.out1(_1956), .in1(R8631), .in2(R8736));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2046 (.out1(_1949), .in1(7 'd 64), .in2(R6295));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2036 (.out1(_1939), .in1(7 'd 64), .in2(R6295));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1992 (.out1(_1898), .in1(R8634), .in2(R8738));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1982 (.out1(_1888), .in1(R8635), .in2(R8739));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1975 (.out1(_1881), .in1(7 'd 64), .in2(R6682));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1964 (.out1(_1870), .in1(R8637), .in2(R8740));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1957 (.out1(_1863), .in1(7 'd 64), .in2(R6682));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1947 (.out1(_1853), .in1(7 'd 64), .in2(R6682));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1903 (.out1(_1812), .in1(R8640), .in2(R8742));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1893 (.out1(_1802), .in1(R8641), .in2(R8743));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1886 (.out1(_1795), .in1(7 'd 64), .in2(R7026));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1875 (.out1(_1784), .in1(R8643), .in2(R8744));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1868 (.out1(_1777), .in1(7 'd 64), .in2(R7026));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1858 (.out1(_1767), .in1(7 'd 64), .in2(R7026));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1814 (.out1(_1726), .in1(R8646), .in2(R8746));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1804 (.out1(_1716), .in1(R8647), .in2(R8747));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1797 (.out1(_1709), .in1(7 'd 64), .in2(R7328));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1786 (.out1(_1698), .in1(R8649), .in2(R8748));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1779 (.out1(_1691), .in1(7 'd 64), .in2(R7328));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1769 (.out1(_1681), .in1(7 'd 64), .in2(R7328));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1725 (.out1(_1640), .in1(R8652), .in2(R8750));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1715 (.out1(_1630), .in1(R8653), .in2(R8751));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1708 (.out1(_1623), .in1(7 'd 64), .in2(R7588));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1697 (.out1(_1612), .in1(R8655), .in2(R8752));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1690 (.out1(_1605), .in1(7 'd 64), .in2(R7588));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1680 (.out1(_1595), .in1(7 'd 64), .in2(R7588));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1636 (.out1(_1554), .in1(R8658), .in2(R8754));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1626 (.out1(_1544), .in1(R8659), .in2(R8755));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1619 (.out1(_1537), .in1(7 'd 64), .in2(R7806));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1608 (.out1(_1526), .in1(R8661), .in2(R8756));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1601 (.out1(_1519), .in1(7 'd 64), .in2(R7806));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1591 (.out1(_1509), .in1(7 'd 64), .in2(R7806));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1547 (.out1(_1468), .in1(R8664), .in2(R8758));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1537 (.out1(_1458), .in1(R8665), .in2(R8759));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1530 (.out1(_1451), .in1(7 'd 64), .in2(R7982));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1519 (.out1(_1440), .in1(R8667), .in2(R8760));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1512 (.out1(_1433), .in1(7 'd 64), .in2(R7982));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1502 (.out1(_1423), .in1(7 'd 64), .in2(R7982));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1458 (.out1(_1382), .in1(R8670), .in2(R8762));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1448 (.out1(_1372), .in1(R8671), .in2(R8763));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1441 (.out1(_1365), .in1(7 'd 64), .in2(R8116));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1430 (.out1(_1354), .in1(R8673), .in2(R8764));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1423 (.out1(_1347), .in1(7 'd 64), .in2(R8116));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1413 (.out1(_1337), .in1(7 'd 64), .in2(R8116));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1369 (.out1(_1296), .in1(R8676), .in2(R8766));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1359 (.out1(_1286), .in1(R8677), .in2(R8767));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1352 (.out1(_1279), .in1(7 'd 64), .in2(R8243));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1341 (.out1(_1268), .in1(R8679), .in2(R8768));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1334 (.out1(_1261), .in1(7 'd 64), .in2(R8243));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1324 (.out1(_1251), .in1(7 'd 64), .in2(R8243));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2562 (.out1(_2447), .in1(b16_bitmap_2528_D), .in2(R8682));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2473 (.out1(_2361), .in1(b24_bitmap_2539_D), .in2(R8683));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2384 (.out1(_2275), .in1(b32_bitmap_2549_D), .in2(R8684));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2295 (.out1(_2189), .in1(b40_bitmap_2559_D), .in2(R8685));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2206 (.out1(_2103), .in1(b48_bitmap_2569_D), .in2(R8686));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2117 (.out1(_2017), .in1(b56_bitmap_2579_D), .in2(R8687));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2089 (.out1(_1992), .in1(_1991), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2000 (.out1(_1906), .in1(_1905), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1911 (.out1(_1820), .in1(_1819), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1822 (.out1(_1734), .in1(_1733), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1733 (.out1(_1648), .in1(_1647), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1644 (.out1(_1562), .in1(_1561), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1555 (.out1(_1476), .in1(_1475), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1466 (.out1(_1390), .in1(_1389), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1377 (.out1(_1304), .in1(_1303), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2621 (.out1(_2506), .in1(R8622), .in2(_2505));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2614 (.out1(_2499), .in1(7 'd 64), .in2(R3081));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2604 (.out1(_2489), .in1(7 'd 64), .in2(R3081));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2586 (.out1(_2471), .in1(7 'd 64), .in2(R3081));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2532 (.out1(_2420), .in1(R8623), .in2(_2419));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2525 (.out1(_2413), .in1(7 'd 64), .in2(R3722));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2515 (.out1(_2403), .in1(7 'd 64), .in2(R3722));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2497 (.out1(_2385), .in1(7 'd 64), .in2(R3722));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2443 (.out1(_2334), .in1(R8624), .in2(_2333));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2436 (.out1(_2327), .in1(7 'd 64), .in2(R4321));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2426 (.out1(_2317), .in1(7 'd 64), .in2(R4321));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2408 (.out1(_2299), .in1(7 'd 64), .in2(R4321));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2354 (.out1(_2248), .in1(R8625), .in2(_2247));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2347 (.out1(_2241), .in1(7 'd 64), .in2(R4878));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2337 (.out1(_2231), .in1(7 'd 64), .in2(R4878));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2319 (.out1(_2213), .in1(7 'd 64), .in2(R4878));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2265 (.out1(_2162), .in1(R8626), .in2(_2161));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2258 (.out1(_2155), .in1(7 'd 64), .in2(R5393));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2248 (.out1(_2145), .in1(7 'd 64), .in2(R5393));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2230 (.out1(_2127), .in1(7 'd 64), .in2(R5393));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2176 (.out1(_2076), .in1(R8627), .in2(_2075));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2169 (.out1(_2069), .in1(7 'd 64), .in2(R5866));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2159 (.out1(_2059), .in1(7 'd 64), .in2(R5866));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2141 (.out1(_2041), .in1(7 'd 64), .in2(R5866));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2090 (.out1(_1993), .in1(_1984), .in2(_1992));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2072 (.out1(_1975), .in1(_1974), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2065 (.out1(_1968), .in1(R8630), .in2(_1967));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2054 (.out1(_1957), .in1(_1956), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2047 (.out1(_1950), .in1(R8632), .in2(_1949));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2037 (.out1(_1940), .in1(R8633), .in2(_1939));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2030 (.out1(_1933), .in1(7 'd 64), .in2(R6295));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2001 (.out1(_1907), .in1(_1898), .in2(_1906));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1983 (.out1(_1889), .in1(_1888), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1976 (.out1(_1882), .in1(R8636), .in2(_1881));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1965 (.out1(_1871), .in1(_1870), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1958 (.out1(_1864), .in1(R8638), .in2(_1863));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1948 (.out1(_1854), .in1(R8639), .in2(_1853));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1941 (.out1(_1847), .in1(7 'd 64), .in2(R6682));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1912 (.out1(_1821), .in1(_1812), .in2(_1820));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1894 (.out1(_1803), .in1(_1802), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1887 (.out1(_1796), .in1(R8642), .in2(_1795));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1876 (.out1(_1785), .in1(_1784), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1869 (.out1(_1778), .in1(R8644), .in2(_1777));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1859 (.out1(_1768), .in1(R8645), .in2(_1767));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1852 (.out1(_1761), .in1(7 'd 64), .in2(R7026));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1823 (.out1(_1735), .in1(_1726), .in2(_1734));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1805 (.out1(_1717), .in1(_1716), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1798 (.out1(_1710), .in1(R8648), .in2(_1709));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1787 (.out1(_1699), .in1(_1698), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1780 (.out1(_1692), .in1(R8650), .in2(_1691));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1770 (.out1(_1682), .in1(R8651), .in2(_1681));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1763 (.out1(_1675), .in1(7 'd 64), .in2(R7328));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1734 (.out1(_1649), .in1(_1640), .in2(_1648));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1716 (.out1(_1631), .in1(_1630), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1709 (.out1(_1624), .in1(R8654), .in2(_1623));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1698 (.out1(_1613), .in1(_1612), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1691 (.out1(_1606), .in1(R8656), .in2(_1605));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1681 (.out1(_1596), .in1(R8657), .in2(_1595));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1674 (.out1(_1589), .in1(7 'd 64), .in2(R7588));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1645 (.out1(_1563), .in1(_1554), .in2(_1562));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1627 (.out1(_1545), .in1(_1544), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1620 (.out1(_1538), .in1(R8660), .in2(_1537));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1609 (.out1(_1527), .in1(_1526), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1602 (.out1(_1520), .in1(R8662), .in2(_1519));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1592 (.out1(_1510), .in1(R8663), .in2(_1509));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1585 (.out1(_1503), .in1(7 'd 64), .in2(R7806));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1556 (.out1(_1477), .in1(_1468), .in2(_1476));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1538 (.out1(_1459), .in1(_1458), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1531 (.out1(_1452), .in1(R8666), .in2(_1451));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1520 (.out1(_1441), .in1(_1440), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1513 (.out1(_1434), .in1(R8668), .in2(_1433));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1503 (.out1(_1424), .in1(R8669), .in2(_1423));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1496 (.out1(_1417), .in1(7 'd 64), .in2(R7982));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1467 (.out1(_1391), .in1(_1382), .in2(_1390));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1449 (.out1(_1373), .in1(_1372), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1442 (.out1(_1366), .in1(R8672), .in2(_1365));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1431 (.out1(_1355), .in1(_1354), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1424 (.out1(_1348), .in1(R8674), .in2(_1347));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1414 (.out1(_1338), .in1(R8675), .in2(_1337));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1407 (.out1(_1331), .in1(7 'd 64), .in2(R8116));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1378 (.out1(_1305), .in1(_1296), .in2(_1304));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1360 (.out1(_1287), .in1(_1286), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1353 (.out1(_1280), .in1(R8678), .in2(_1279));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1342 (.out1(_1269), .in1(_1268), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1335 (.out1(_1262), .in1(R8680), .in2(_1261));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1325 (.out1(_1252), .in1(R8681), .in2(_1251));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1318 (.out1(_1245), .in1(7 'd 64), .in2(R8243));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2875 (.out1(R2876), .clock(clock), .in1(R2875));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3081 (.out1(R3082), .clock(clock), .in1(R3081));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3283 (.out1(R3284), .clock(clock), .in1(R3283));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3530 (.out1(R3531), .clock(clock), .in1(R3530));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3722 (.out1(R3723), .clock(clock), .in1(R3722));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3910 (.out1(R3911), .clock(clock), .in1(R3910));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4143 (.out1(R4144), .clock(clock), .in1(R4143));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4321 (.out1(R4322), .clock(clock), .in1(R4321));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4495 (.out1(R4496), .clock(clock), .in1(R4495));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4714 (.out1(R4715), .clock(clock), .in1(R4714));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4878 (.out1(R4879), .clock(clock), .in1(R4878));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5038 (.out1(R5039), .clock(clock), .in1(R5038));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5243 (.out1(R5244), .clock(clock), .in1(R5243));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5393 (.out1(R5394), .clock(clock), .in1(R5393));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5539 (.out1(R5540), .clock(clock), .in1(R5539));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5730 (.out1(R5731), .clock(clock), .in1(R5730));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5866 (.out1(R5867), .clock(clock), .in1(R5866));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5998 (.out1(R5999), .clock(clock), .in1(R5998));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6174 (.out1(R6175), .clock(clock), .in1(R6174));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6412 (.out1(R6413), .clock(clock), .in1(R6412));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6575 (.out1(R6576), .clock(clock), .in1(R6575));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6785 (.out1(R6786), .clock(clock), .in1(R6785));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6933 (.out1(R6934), .clock(clock), .in1(R6933));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7115 (.out1(R7116), .clock(clock), .in1(R7115));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7249 (.out1(R7250), .clock(clock), .in1(R7249));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7403 (.out1(R7404), .clock(clock), .in1(R7403));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7523 (.out1(R7524), .clock(clock), .in1(R7523));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7649 (.out1(R7650), .clock(clock), .in1(R7649));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7755 (.out1(R7756), .clock(clock), .in1(R7755));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7853 (.out1(R7854), .clock(clock), .in1(R7853));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7945 (.out1(R7946), .clock(clock), .in1(R7945));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8015 (.out1(R8016), .clock(clock), .in1(R8015));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8093 (.out1(R8094), .clock(clock), .in1(R8093));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8135 (.out1(R8136), .clock(clock), .in1(R8135));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8198 (.out1(R8199), .clock(clock), .in1(R8198));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8262 (.out1(R8263), .clock(clock), .in1(R8262));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8273 (.out1(R8274), .clock(clock), .in1(R8273));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8284 (.out1(R8285), .clock(clock), .in1(R8284));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8295 (.out1(R8296), .clock(clock), .in1(R8295));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8306 (.out1(R8307), .clock(clock), .in1(R8306));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8317 (.out1(R8318), .clock(clock), .in1(R8317));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8328 (.out1(R8329), .clock(clock), .in1(R8328));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8339 (.out1(R8340), .clock(clock), .in1(R8339));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8350 (.out1(R8351), .clock(clock), .in1(R8350));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8375 (.out1(R8376), .clock(clock), .in1(R8375));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8386 (.out1(R8387), .clock(clock), .in1(R8386));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8397 (.out1(R8398), .clock(clock), .in1(R8397));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8408 (.out1(R8409), .clock(clock), .in1(R8408));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8419 (.out1(R8420), .clock(clock), .in1(R8419));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8430 (.out1(R8431), .clock(clock), .in1(R8430));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8768 (.out1(R8769), .clock(clock), .in1(_2498));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8769 (.out1(R8770), .clock(clock), .in1(_2488));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8770 (.out1(R8771), .clock(clock), .in1(_2482));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8771 (.out1(R8772), .clock(clock), .in1(_2470));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8772 (.out1(R8773), .clock(clock), .in1(_2464));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8773 (.out1(R8774), .clock(clock), .in1(_2454));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8774 (.out1(R8775), .clock(clock), .in1(_2412));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8775 (.out1(R8776), .clock(clock), .in1(_2402));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8776 (.out1(R8777), .clock(clock), .in1(_2396));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8777 (.out1(R8778), .clock(clock), .in1(_2384));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8778 (.out1(R8779), .clock(clock), .in1(_2378));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8779 (.out1(R8780), .clock(clock), .in1(_2368));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8780 (.out1(R8781), .clock(clock), .in1(_2326));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8781 (.out1(R8782), .clock(clock), .in1(_2316));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8782 (.out1(R8783), .clock(clock), .in1(_2310));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8783 (.out1(R8784), .clock(clock), .in1(_2298));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8784 (.out1(R8785), .clock(clock), .in1(_2292));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8785 (.out1(R8786), .clock(clock), .in1(_2282));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8786 (.out1(R8787), .clock(clock), .in1(_2240));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8787 (.out1(R8788), .clock(clock), .in1(_2230));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8788 (.out1(R8789), .clock(clock), .in1(_2224));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8789 (.out1(R8790), .clock(clock), .in1(_2212));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8790 (.out1(R8791), .clock(clock), .in1(_2206));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8791 (.out1(R8792), .clock(clock), .in1(_2196));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8792 (.out1(R8793), .clock(clock), .in1(_2154));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8793 (.out1(R8794), .clock(clock), .in1(_2144));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8794 (.out1(R8795), .clock(clock), .in1(_2138));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8795 (.out1(R8796), .clock(clock), .in1(_2126));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8796 (.out1(R8797), .clock(clock), .in1(_2120));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8797 (.out1(R8798), .clock(clock), .in1(_2110));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8798 (.out1(R8799), .clock(clock), .in1(_2068));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8799 (.out1(R8800), .clock(clock), .in1(_2058));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8800 (.out1(R8801), .clock(clock), .in1(_2052));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8801 (.out1(R8802), .clock(clock), .in1(_2040));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8802 (.out1(R8803), .clock(clock), .in1(_2034));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8803 (.out1(R8804), .clock(clock), .in1(_2024));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8804 (.out1(R8805), .clock(clock), .in1(_1932));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8805 (.out1(R8806), .clock(clock), .in1(_1846));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8806 (.out1(R8807), .clock(clock), .in1(_1760));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8807 (.out1(R8808), .clock(clock), .in1(_1674));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8808 (.out1(R8809), .clock(clock), .in1(_1588));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8809 (.out1(R8810), .clock(clock), .in1(_1502));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8810 (.out1(R8811), .clock(clock), .in1(_1416));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8811 (.out1(R8812), .clock(clock), .in1(_1330));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8812 (.out1(R8813), .clock(clock), .in1(_1244));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8813 (.out1(R8814), .clock(clock), .in1(_2447));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8814 (.out1(R8815), .clock(clock), .in1(_2361));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8815 (.out1(R8816), .clock(clock), .in1(_2275));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8816 (.out1(R8817), .clock(clock), .in1(_2189));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8817 (.out1(R8818), .clock(clock), .in1(_2103));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8818 (.out1(R8819), .clock(clock), .in1(_2017));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8819 (.out1(R8820), .clock(clock), .in1(_2506));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8820 (.out1(R8821), .clock(clock), .in1(_2499));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8821 (.out1(R8822), .clock(clock), .in1(_2489));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8822 (.out1(R8823), .clock(clock), .in1(_2471));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8823 (.out1(R8824), .clock(clock), .in1(_2420));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8824 (.out1(R8825), .clock(clock), .in1(_2413));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8825 (.out1(R8826), .clock(clock), .in1(_2403));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8826 (.out1(R8827), .clock(clock), .in1(_2385));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8827 (.out1(R8828), .clock(clock), .in1(_2334));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8828 (.out1(R8829), .clock(clock), .in1(_2327));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8829 (.out1(R8830), .clock(clock), .in1(_2317));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8830 (.out1(R8831), .clock(clock), .in1(_2299));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8831 (.out1(R8832), .clock(clock), .in1(_2248));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8832 (.out1(R8833), .clock(clock), .in1(_2241));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8833 (.out1(R8834), .clock(clock), .in1(_2231));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8834 (.out1(R8835), .clock(clock), .in1(_2213));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8835 (.out1(R8836), .clock(clock), .in1(_2162));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8836 (.out1(R8837), .clock(clock), .in1(_2155));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8837 (.out1(R8838), .clock(clock), .in1(_2145));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8838 (.out1(R8839), .clock(clock), .in1(_2127));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8839 (.out1(R8840), .clock(clock), .in1(_2076));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8840 (.out1(R8841), .clock(clock), .in1(_2069));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8841 (.out1(R8842), .clock(clock), .in1(_2059));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8842 (.out1(R8843), .clock(clock), .in1(_2041));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8843 (.out1(R8844), .clock(clock), .in1(_1993));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8844 (.out1(R8845), .clock(clock), .in1(_1975));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8845 (.out1(R8846), .clock(clock), .in1(_1968));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8846 (.out1(R8847), .clock(clock), .in1(_1957));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8847 (.out1(R8848), .clock(clock), .in1(_1950));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8848 (.out1(R8849), .clock(clock), .in1(_1940));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8849 (.out1(R8850), .clock(clock), .in1(_1933));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8850 (.out1(R8851), .clock(clock), .in1(_1907));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8851 (.out1(R8852), .clock(clock), .in1(_1889));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8852 (.out1(R8853), .clock(clock), .in1(_1882));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8853 (.out1(R8854), .clock(clock), .in1(_1871));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8854 (.out1(R8855), .clock(clock), .in1(_1864));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8855 (.out1(R8856), .clock(clock), .in1(_1854));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8856 (.out1(R8857), .clock(clock), .in1(_1847));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8857 (.out1(R8858), .clock(clock), .in1(_1821));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8858 (.out1(R8859), .clock(clock), .in1(_1803));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8859 (.out1(R8860), .clock(clock), .in1(_1796));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8860 (.out1(R8861), .clock(clock), .in1(_1785));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8861 (.out1(R8862), .clock(clock), .in1(_1778));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8862 (.out1(R8863), .clock(clock), .in1(_1768));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8863 (.out1(R8864), .clock(clock), .in1(_1761));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8864 (.out1(R8865), .clock(clock), .in1(_1735));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8865 (.out1(R8866), .clock(clock), .in1(_1717));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8866 (.out1(R8867), .clock(clock), .in1(_1710));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8867 (.out1(R8868), .clock(clock), .in1(_1699));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8868 (.out1(R8869), .clock(clock), .in1(_1692));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8869 (.out1(R8870), .clock(clock), .in1(_1682));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8870 (.out1(R8871), .clock(clock), .in1(_1675));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8871 (.out1(R8872), .clock(clock), .in1(_1649));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8872 (.out1(R8873), .clock(clock), .in1(_1631));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8873 (.out1(R8874), .clock(clock), .in1(_1624));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8874 (.out1(R8875), .clock(clock), .in1(_1613));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8875 (.out1(R8876), .clock(clock), .in1(_1606));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8876 (.out1(R8877), .clock(clock), .in1(_1596));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8877 (.out1(R8878), .clock(clock), .in1(_1589));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8878 (.out1(R8879), .clock(clock), .in1(_1563));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8879 (.out1(R8880), .clock(clock), .in1(_1545));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8880 (.out1(R8881), .clock(clock), .in1(_1538));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8881 (.out1(R8882), .clock(clock), .in1(_1527));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8882 (.out1(R8883), .clock(clock), .in1(_1520));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8883 (.out1(R8884), .clock(clock), .in1(_1510));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8884 (.out1(R8885), .clock(clock), .in1(_1503));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8885 (.out1(R8886), .clock(clock), .in1(_1477));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8886 (.out1(R8887), .clock(clock), .in1(_1459));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8887 (.out1(R8888), .clock(clock), .in1(_1452));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8888 (.out1(R8889), .clock(clock), .in1(_1441));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8889 (.out1(R8890), .clock(clock), .in1(_1434));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8890 (.out1(R8891), .clock(clock), .in1(_1424));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8891 (.out1(R8892), .clock(clock), .in1(_1417));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8892 (.out1(R8893), .clock(clock), .in1(_1391));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8893 (.out1(R8894), .clock(clock), .in1(_1373));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8894 (.out1(R8895), .clock(clock), .in1(_1366));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8895 (.out1(R8896), .clock(clock), .in1(_1355));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8896 (.out1(R8897), .clock(clock), .in1(_1348));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8897 (.out1(R8898), .clock(clock), .in1(_1338));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8898 (.out1(R8899), .clock(clock), .in1(_1331));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8899 (.out1(R8900), .clock(clock), .in1(_1305));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8900 (.out1(R8901), .clock(clock), .in1(_1287));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8901 (.out1(R8902), .clock(clock), .in1(_1280));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8902 (.out1(R8903), .clock(clock), .in1(_1269));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8903 (.out1(R8904), .clock(clock), .in1(_1262));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8904 (.out1(R8905), .clock(clock), .in1(_1252));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8905 (.out1(R8906), .clock(clock), .in1(_1245));
  SRAM op2563 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2448),.ADR(R8814));
  SRAM op2474 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2362),.ADR(R8815));
  SRAM op2385 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2276),.ADR(R8816));
  SRAM op2296 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2190),.ADR(R8817));
  SRAM op2207 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2104),.ADR(R8818));
  SRAM op2118 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2018),.ADR(R8819));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2022 (.out1(_1925), .in1(R6175));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1933 (.out1(_1839), .in1(R6576));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1844 (.out1(_1753), .in1(R6934));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1755 (.out1(_1667), .in1(R7250));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1666 (.out1(_1581), .in1(R7524));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1577 (.out1(_1495), .in1(R7756));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1488 (.out1(_1409), .in1(R7946));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1399 (.out1(_1323), .in1(R8094));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1310 (.out1(_1237), .in1(R8199));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2073 (.out1(_1976), .in1(R8845), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1984 (.out1(_1890), .in1(R8852), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1895 (.out1(_1804), .in1(R8859), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1806 (.out1(_1718), .in1(R8866), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1717 (.out1(_1632), .in1(R8873), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1628 (.out1(_1546), .in1(R8880), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1539 (.out1(_1460), .in1(R8887), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1450 (.out1(_1374), .in1(R8894), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1361 (.out1(_1288), .in1(R8901), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2622 (.out1(_2507), .in1(R8820), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2533 (.out1(_2421), .in1(R8824), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2444 (.out1(_2335), .in1(R8828), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2355 (.out1(_2249), .in1(R8832), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2266 (.out1(_2163), .in1(R8836), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2177 (.out1(_2077), .in1(R8840), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2091 (.out1(_1994), .in1(R8844), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2074 (.out1(_1977), .in1(R8846), .in2(_1976));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2055 (.out1(_1958), .in1(R8847), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2038 (.out1(_1941), .in1(R8849), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2002 (.out1(_1908), .in1(R8851), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1985 (.out1(_1891), .in1(R8853), .in2(_1890));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1966 (.out1(_1872), .in1(R8854), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1949 (.out1(_1855), .in1(R8856), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1913 (.out1(_1822), .in1(R8858), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1896 (.out1(_1805), .in1(R8860), .in2(_1804));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1877 (.out1(_1786), .in1(R8861), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1860 (.out1(_1769), .in1(R8863), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1824 (.out1(_1736), .in1(R8865), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1807 (.out1(_1719), .in1(R8867), .in2(_1718));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1788 (.out1(_1700), .in1(R8868), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1771 (.out1(_1683), .in1(R8870), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1735 (.out1(_1650), .in1(R8872), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1718 (.out1(_1633), .in1(R8874), .in2(_1632));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1699 (.out1(_1614), .in1(R8875), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1682 (.out1(_1597), .in1(R8877), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1646 (.out1(_1564), .in1(R8879), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1629 (.out1(_1547), .in1(R8881), .in2(_1546));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1610 (.out1(_1528), .in1(R8882), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1593 (.out1(_1511), .in1(R8884), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1557 (.out1(_1478), .in1(R8886), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1540 (.out1(_1461), .in1(R8888), .in2(_1460));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1521 (.out1(_1442), .in1(R8889), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1504 (.out1(_1425), .in1(R8891), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1468 (.out1(_1392), .in1(R8893), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1451 (.out1(_1375), .in1(R8895), .in2(_1374));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1432 (.out1(_1356), .in1(R8896), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1415 (.out1(_1339), .in1(R8898), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1379 (.out1(_1306), .in1(R8900), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1362 (.out1(_1289), .in1(R8902), .in2(_1288));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1343 (.out1(_1270), .in1(R8903), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1326 (.out1(_1253), .in1(R8905), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2615 (.out1(_2500), .in1(R8769), .in2(R8821));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2605 (.out1(_2490), .in1(R8770), .in2(R8822));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2598 (.out1(_2483), .in1(7 'd 64), .in2(R3082));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2587 (.out1(_2472), .in1(R8772), .in2(R8823));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2580 (.out1(_2465), .in1(7 'd 64), .in2(R3082));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2570 (.out1(_2455), .in1(7 'd 64), .in2(R3082));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2526 (.out1(_2414), .in1(R8775), .in2(R8825));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2516 (.out1(_2404), .in1(R8776), .in2(R8826));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2509 (.out1(_2397), .in1(7 'd 64), .in2(R3723));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2498 (.out1(_2386), .in1(R8778), .in2(R8827));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2491 (.out1(_2379), .in1(7 'd 64), .in2(R3723));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2481 (.out1(_2369), .in1(7 'd 64), .in2(R3723));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2437 (.out1(_2328), .in1(R8781), .in2(R8829));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2427 (.out1(_2318), .in1(R8782), .in2(R8830));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2420 (.out1(_2311), .in1(7 'd 64), .in2(R4322));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2409 (.out1(_2300), .in1(R8784), .in2(R8831));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2402 (.out1(_2293), .in1(7 'd 64), .in2(R4322));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2392 (.out1(_2283), .in1(7 'd 64), .in2(R4322));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2348 (.out1(_2242), .in1(R8787), .in2(R8833));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2338 (.out1(_2232), .in1(R8788), .in2(R8834));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2331 (.out1(_2225), .in1(7 'd 64), .in2(R4879));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2320 (.out1(_2214), .in1(R8790), .in2(R8835));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2313 (.out1(_2207), .in1(7 'd 64), .in2(R4879));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2303 (.out1(_2197), .in1(7 'd 64), .in2(R4879));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2259 (.out1(_2156), .in1(R8793), .in2(R8837));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2249 (.out1(_2146), .in1(R8794), .in2(R8838));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2242 (.out1(_2139), .in1(7 'd 64), .in2(R5394));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2231 (.out1(_2128), .in1(R8796), .in2(R8839));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2224 (.out1(_2121), .in1(7 'd 64), .in2(R5394));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2214 (.out1(_2111), .in1(7 'd 64), .in2(R5394));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2170 (.out1(_2070), .in1(R8799), .in2(R8841));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2160 (.out1(_2060), .in1(R8800), .in2(R8842));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2153 (.out1(_2053), .in1(7 'd 64), .in2(R5867));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2142 (.out1(_2042), .in1(R8802), .in2(R8843));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2135 (.out1(_2035), .in1(7 'd 64), .in2(R5867));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2125 (.out1(_2025), .in1(7 'd 64), .in2(R5867));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2056 (.out1(_1959), .in1(R8848), .in2(_1958));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2031 (.out1(_1934), .in1(R8805), .in2(R8850));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1967 (.out1(_1873), .in1(R8855), .in2(_1872));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1942 (.out1(_1848), .in1(R8806), .in2(R8857));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1878 (.out1(_1787), .in1(R8862), .in2(_1786));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1853 (.out1(_1762), .in1(R8807), .in2(R8864));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1789 (.out1(_1701), .in1(R8869), .in2(_1700));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1764 (.out1(_1676), .in1(R8808), .in2(R8871));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1700 (.out1(_1615), .in1(R8876), .in2(_1614));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1675 (.out1(_1590), .in1(R8809), .in2(R8878));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1611 (.out1(_1529), .in1(R8883), .in2(_1528));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1586 (.out1(_1504), .in1(R8810), .in2(R8885));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1522 (.out1(_1443), .in1(R8890), .in2(_1442));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1497 (.out1(_1418), .in1(R8811), .in2(R8892));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1433 (.out1(_1357), .in1(R8897), .in2(_1356));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1408 (.out1(_1332), .in1(R8812), .in2(R8899));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1344 (.out1(_1271), .in1(R8904), .in2(_1270));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1319 (.out1(_1246), .in1(R8813), .in2(R8906));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2023 (.out1(_1926), .in1(_1925), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1934 (.out1(_1840), .in1(_1839), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1845 (.out1(_1754), .in1(_1753), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1756 (.out1(_1668), .in1(_1667), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1667 (.out1(_1582), .in1(_1581), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1578 (.out1(_1496), .in1(_1495), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1489 (.out1(_1410), .in1(_1409), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1400 (.out1(_1324), .in1(_1323), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1311 (.out1(_1238), .in1(_1237), .in2(2 'd 2));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2623 (.out1(_2508), .in1(_2507), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2534 (.out1(_2422), .in1(_2421), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2445 (.out1(_2336), .in1(_2335), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2356 (.out1(_2250), .in1(_2249), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2267 (.out1(_2164), .in1(_2163), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2178 (.out1(_2078), .in1(_2077), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2092 (.out1(_1995), .in1(_1994), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2075 (.out1(_1978), .in1(_1977), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2039 (.out1(_1942), .in1(_1941), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2003 (.out1(_1909), .in1(_1908), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1986 (.out1(_1892), .in1(_1891), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1950 (.out1(_1856), .in1(_1855), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1914 (.out1(_1823), .in1(_1822), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1897 (.out1(_1806), .in1(_1805), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1861 (.out1(_1770), .in1(_1769), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1825 (.out1(_1737), .in1(_1736), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1808 (.out1(_1720), .in1(_1719), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1772 (.out1(_1684), .in1(_1683), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1736 (.out1(_1651), .in1(_1650), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1719 (.out1(_1634), .in1(_1633), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1683 (.out1(_1598), .in1(_1597), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1647 (.out1(_1565), .in1(_1564), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1630 (.out1(_1548), .in1(_1547), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1594 (.out1(_1512), .in1(_1511), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1558 (.out1(_1479), .in1(_1478), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1541 (.out1(_1462), .in1(_1461), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1505 (.out1(_1426), .in1(_1425), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1469 (.out1(_1393), .in1(_1392), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1452 (.out1(_1376), .in1(_1375), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1416 (.out1(_1340), .in1(_1339), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1380 (.out1(_1307), .in1(_1306), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1363 (.out1(_1290), .in1(_1289), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1327 (.out1(_1254), .in1(_1253), .in2(63 'd 6148914691236517205));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2624 (.out1(_2509), .in1(_2500), .in2(_2508));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2606 (.out1(_2491), .in1(_2490), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2599 (.out1(_2484), .in1(R8771), .in2(_2483));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2588 (.out1(_2473), .in1(_2472), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2581 (.out1(_2466), .in1(R8773), .in2(_2465));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2571 (.out1(_2456), .in1(R8774), .in2(_2455));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2564 (.out1(_2449), .in1(7 'd 64), .in2(R3082));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2535 (.out1(_2423), .in1(_2414), .in2(_2422));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2517 (.out1(_2405), .in1(_2404), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2510 (.out1(_2398), .in1(R8777), .in2(_2397));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2499 (.out1(_2387), .in1(_2386), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2492 (.out1(_2380), .in1(R8779), .in2(_2379));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2482 (.out1(_2370), .in1(R8780), .in2(_2369));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2475 (.out1(_2363), .in1(7 'd 64), .in2(R3723));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2446 (.out1(_2337), .in1(_2328), .in2(_2336));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2428 (.out1(_2319), .in1(_2318), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2421 (.out1(_2312), .in1(R8783), .in2(_2311));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2410 (.out1(_2301), .in1(_2300), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2403 (.out1(_2294), .in1(R8785), .in2(_2293));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2393 (.out1(_2284), .in1(R8786), .in2(_2283));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2386 (.out1(_2277), .in1(7 'd 64), .in2(R4322));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2357 (.out1(_2251), .in1(_2242), .in2(_2250));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2339 (.out1(_2233), .in1(_2232), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2332 (.out1(_2226), .in1(R8789), .in2(_2225));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2321 (.out1(_2215), .in1(_2214), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2314 (.out1(_2208), .in1(R8791), .in2(_2207));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2304 (.out1(_2198), .in1(R8792), .in2(_2197));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2297 (.out1(_2191), .in1(7 'd 64), .in2(R4879));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2268 (.out1(_2165), .in1(_2156), .in2(_2164));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2250 (.out1(_2147), .in1(_2146), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2243 (.out1(_2140), .in1(R8795), .in2(_2139));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2232 (.out1(_2129), .in1(_2128), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2225 (.out1(_2122), .in1(R8797), .in2(_2121));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2215 (.out1(_2112), .in1(R8798), .in2(_2111));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2208 (.out1(_2105), .in1(7 'd 64), .in2(R5394));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2179 (.out1(_2079), .in1(_2070), .in2(_2078));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2161 (.out1(_2061), .in1(_2060), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2154 (.out1(_2054), .in1(R8801), .in2(_2053));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2143 (.out1(_2043), .in1(_2042), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2136 (.out1(_2036), .in1(R8803), .in2(_2035));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2126 (.out1(_2026), .in1(R8804), .in2(_2025));
  SUB_GATE #(.BITSIZE_in1(7), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2119 (.out1(_2019), .in1(7 'd 64), .in2(R5867));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2093 (.out1(_1996), .in1(_1978), .in2(_1995));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2057 (.out1(_1960), .in1(_1959), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2040 (.out1(_1943), .in1(_1934), .in2(_1942));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2004 (.out1(_1910), .in1(_1892), .in2(_1909));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1968 (.out1(_1874), .in1(_1873), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1951 (.out1(_1857), .in1(_1848), .in2(_1856));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1915 (.out1(_1824), .in1(_1806), .in2(_1823));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1879 (.out1(_1788), .in1(_1787), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1862 (.out1(_1771), .in1(_1762), .in2(_1770));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1826 (.out1(_1738), .in1(_1720), .in2(_1737));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1790 (.out1(_1702), .in1(_1701), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1773 (.out1(_1685), .in1(_1676), .in2(_1684));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1737 (.out1(_1652), .in1(_1634), .in2(_1651));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1701 (.out1(_1616), .in1(_1615), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1684 (.out1(_1599), .in1(_1590), .in2(_1598));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1648 (.out1(_1566), .in1(_1548), .in2(_1565));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1612 (.out1(_1530), .in1(_1529), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1595 (.out1(_1513), .in1(_1504), .in2(_1512));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1559 (.out1(_1480), .in1(_1462), .in2(_1479));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1523 (.out1(_1444), .in1(_1443), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1506 (.out1(_1427), .in1(_1418), .in2(_1426));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1470 (.out1(_1394), .in1(_1376), .in2(_1393));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1434 (.out1(_1358), .in1(_1357), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1417 (.out1(_1341), .in1(_1332), .in2(_1340));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1381 (.out1(_1308), .in1(_1290), .in2(_1307));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1345 (.out1(_1272), .in1(_1271), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1328 (.out1(_1255), .in1(_1246), .in2(_1254));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op2876 (.out1(R2877), .clock(clock), .in1(R2876));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3284 (.out1(R3285), .clock(clock), .in1(R3284));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3531 (.out1(R3532), .clock(clock), .in1(R3531));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3911 (.out1(R3912), .clock(clock), .in1(R3911));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4144 (.out1(R4145), .clock(clock), .in1(R4144));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4496 (.out1(R4497), .clock(clock), .in1(R4496));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4715 (.out1(R4716), .clock(clock), .in1(R4715));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5039 (.out1(R5040), .clock(clock), .in1(R5039));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5244 (.out1(R5245), .clock(clock), .in1(R5244));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5540 (.out1(R5541), .clock(clock), .in1(R5540));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5731 (.out1(R5732), .clock(clock), .in1(R5731));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5999 (.out1(R6000), .clock(clock), .in1(R5999));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6413 (.out1(R6414), .clock(clock), .in1(R6413));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6786 (.out1(R6787), .clock(clock), .in1(R6786));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7116 (.out1(R7117), .clock(clock), .in1(R7116));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7404 (.out1(R7405), .clock(clock), .in1(R7404));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7650 (.out1(R7651), .clock(clock), .in1(R7650));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7854 (.out1(R7855), .clock(clock), .in1(R7854));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8016 (.out1(R8017), .clock(clock), .in1(R8016));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8136 (.out1(R8137), .clock(clock), .in1(R8136));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8263 (.out1(R8264), .clock(clock), .in1(R8263));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8274 (.out1(R8275), .clock(clock), .in1(R8274));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8285 (.out1(R8286), .clock(clock), .in1(R8285));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8296 (.out1(R8297), .clock(clock), .in1(R8296));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8307 (.out1(R8308), .clock(clock), .in1(R8307));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8318 (.out1(R8319), .clock(clock), .in1(R8318));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8329 (.out1(R8330), .clock(clock), .in1(R8329));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8340 (.out1(R8341), .clock(clock), .in1(R8340));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8351 (.out1(R8352), .clock(clock), .in1(R8351));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8376 (.out1(R8377), .clock(clock), .in1(R8376));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8387 (.out1(R8388), .clock(clock), .in1(R8387));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8398 (.out1(R8399), .clock(clock), .in1(R8398));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8409 (.out1(R8410), .clock(clock), .in1(R8409));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8420 (.out1(R8421), .clock(clock), .in1(R8420));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8431 (.out1(R8432), .clock(clock), .in1(R8431));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8906 (.out1(R8907), .clock(clock), .in1(_2448));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8907 (.out1(R8908), .clock(clock), .in1(_2362));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8908 (.out1(R8909), .clock(clock), .in1(_2276));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8909 (.out1(R8910), .clock(clock), .in1(_2190));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8910 (.out1(R8911), .clock(clock), .in1(_2104));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8911 (.out1(R8912), .clock(clock), .in1(_2018));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8912 (.out1(R8913), .clock(clock), .in1(_1926));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8913 (.out1(R8914), .clock(clock), .in1(_1840));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8914 (.out1(R8915), .clock(clock), .in1(_1754));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8915 (.out1(R8916), .clock(clock), .in1(_1668));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8916 (.out1(R8917), .clock(clock), .in1(_1582));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8917 (.out1(R8918), .clock(clock), .in1(_1496));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8918 (.out1(R8919), .clock(clock), .in1(_1410));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8919 (.out1(R8920), .clock(clock), .in1(_1324));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8920 (.out1(R8921), .clock(clock), .in1(_1238));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8921 (.out1(R8922), .clock(clock), .in1(_2509));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8922 (.out1(R8923), .clock(clock), .in1(_2491));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8923 (.out1(R8924), .clock(clock), .in1(_2484));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8924 (.out1(R8925), .clock(clock), .in1(_2473));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8925 (.out1(R8926), .clock(clock), .in1(_2466));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8926 (.out1(R8927), .clock(clock), .in1(_2456));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8927 (.out1(R8928), .clock(clock), .in1(_2449));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8928 (.out1(R8929), .clock(clock), .in1(_2423));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8929 (.out1(R8930), .clock(clock), .in1(_2405));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8930 (.out1(R8931), .clock(clock), .in1(_2398));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8931 (.out1(R8932), .clock(clock), .in1(_2387));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8932 (.out1(R8933), .clock(clock), .in1(_2380));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8933 (.out1(R8934), .clock(clock), .in1(_2370));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8934 (.out1(R8935), .clock(clock), .in1(_2363));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8935 (.out1(R8936), .clock(clock), .in1(_2337));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8936 (.out1(R8937), .clock(clock), .in1(_2319));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8937 (.out1(R8938), .clock(clock), .in1(_2312));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8938 (.out1(R8939), .clock(clock), .in1(_2301));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8939 (.out1(R8940), .clock(clock), .in1(_2294));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8940 (.out1(R8941), .clock(clock), .in1(_2284));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8941 (.out1(R8942), .clock(clock), .in1(_2277));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8942 (.out1(R8943), .clock(clock), .in1(_2251));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8943 (.out1(R8944), .clock(clock), .in1(_2233));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8944 (.out1(R8945), .clock(clock), .in1(_2226));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8945 (.out1(R8946), .clock(clock), .in1(_2215));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8946 (.out1(R8947), .clock(clock), .in1(_2208));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8947 (.out1(R8948), .clock(clock), .in1(_2198));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8948 (.out1(R8949), .clock(clock), .in1(_2191));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8949 (.out1(R8950), .clock(clock), .in1(_2165));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8950 (.out1(R8951), .clock(clock), .in1(_2147));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8951 (.out1(R8952), .clock(clock), .in1(_2140));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8952 (.out1(R8953), .clock(clock), .in1(_2129));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8953 (.out1(R8954), .clock(clock), .in1(_2122));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8954 (.out1(R8955), .clock(clock), .in1(_2112));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8955 (.out1(R8956), .clock(clock), .in1(_2105));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8956 (.out1(R8957), .clock(clock), .in1(_2079));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8957 (.out1(R8958), .clock(clock), .in1(_2061));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8958 (.out1(R8959), .clock(clock), .in1(_2054));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8959 (.out1(R8960), .clock(clock), .in1(_2043));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8960 (.out1(R8961), .clock(clock), .in1(_2036));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8961 (.out1(R8962), .clock(clock), .in1(_2026));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8962 (.out1(R8963), .clock(clock), .in1(_2019));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8963 (.out1(R8964), .clock(clock), .in1(_1996));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8964 (.out1(R8965), .clock(clock), .in1(_1960));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8965 (.out1(R8966), .clock(clock), .in1(_1943));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8966 (.out1(R8967), .clock(clock), .in1(_1910));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8967 (.out1(R8968), .clock(clock), .in1(_1874));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8968 (.out1(R8969), .clock(clock), .in1(_1857));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8969 (.out1(R8970), .clock(clock), .in1(_1824));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8970 (.out1(R8971), .clock(clock), .in1(_1788));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8971 (.out1(R8972), .clock(clock), .in1(_1771));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8972 (.out1(R8973), .clock(clock), .in1(_1738));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8973 (.out1(R8974), .clock(clock), .in1(_1702));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8974 (.out1(R8975), .clock(clock), .in1(_1685));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8975 (.out1(R8976), .clock(clock), .in1(_1652));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8976 (.out1(R8977), .clock(clock), .in1(_1616));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8977 (.out1(R8978), .clock(clock), .in1(_1599));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8978 (.out1(R8979), .clock(clock), .in1(_1566));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8979 (.out1(R8980), .clock(clock), .in1(_1530));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8980 (.out1(R8981), .clock(clock), .in1(_1513));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8981 (.out1(R8982), .clock(clock), .in1(_1480));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8982 (.out1(R8983), .clock(clock), .in1(_1444));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8983 (.out1(R8984), .clock(clock), .in1(_1427));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8984 (.out1(R8985), .clock(clock), .in1(_1394));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8985 (.out1(R8986), .clock(clock), .in1(_1358));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8986 (.out1(R8987), .clock(clock), .in1(_1341));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8987 (.out1(R8988), .clock(clock), .in1(_1308));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8988 (.out1(R8989), .clock(clock), .in1(_1272));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8989 (.out1(R8990), .clock(clock), .in1(_1255));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2556 (.out1(_2441), .in1(R2877));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2467 (.out1(_2355), .in1(R3532));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2378 (.out1(_2269), .in1(R4145));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2289 (.out1(_2183), .in1(R4716));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2200 (.out1(_2097), .in1(R5245));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2111 (.out1(_2011), .in1(R5732));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2607 (.out1(_2492), .in1(R8923), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2518 (.out1(_2406), .in1(R8930), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2429 (.out1(_2320), .in1(R8937), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2340 (.out1(_2234), .in1(R8944), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2251 (.out1(_2148), .in1(R8951), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2162 (.out1(_2062), .in1(R8958), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2058 (.out1(_1961), .in1(R8965), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2041 (.out1(_1944), .in1(R8966), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1969 (.out1(_1875), .in1(R8968), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1952 (.out1(_1858), .in1(R8969), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1880 (.out1(_1789), .in1(R8971), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1863 (.out1(_1772), .in1(R8972), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1791 (.out1(_1703), .in1(R8974), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1774 (.out1(_1686), .in1(R8975), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1702 (.out1(_1617), .in1(R8977), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1685 (.out1(_1600), .in1(R8978), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1613 (.out1(_1531), .in1(R8980), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1596 (.out1(_1514), .in1(R8981), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1524 (.out1(_1445), .in1(R8983), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1507 (.out1(_1428), .in1(R8984), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1435 (.out1(_1359), .in1(R8986), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1418 (.out1(_1342), .in1(R8987), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1346 (.out1(_1273), .in1(R8989), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1329 (.out1(_1256), .in1(R8990), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2625 (.out1(_2510), .in1(R8922), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2608 (.out1(_2493), .in1(R8924), .in2(_2492));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2589 (.out1(_2474), .in1(R8925), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2572 (.out1(_2457), .in1(R8927), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2536 (.out1(_2424), .in1(R8929), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2519 (.out1(_2407), .in1(R8931), .in2(_2406));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2500 (.out1(_2388), .in1(R8932), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2483 (.out1(_2371), .in1(R8934), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2447 (.out1(_2338), .in1(R8936), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2430 (.out1(_2321), .in1(R8938), .in2(_2320));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2411 (.out1(_2302), .in1(R8939), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2394 (.out1(_2285), .in1(R8941), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2358 (.out1(_2252), .in1(R8943), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2341 (.out1(_2235), .in1(R8945), .in2(_2234));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2322 (.out1(_2216), .in1(R8946), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2305 (.out1(_2199), .in1(R8948), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2269 (.out1(_2166), .in1(R8950), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2252 (.out1(_2149), .in1(R8952), .in2(_2148));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2233 (.out1(_2130), .in1(R8953), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2216 (.out1(_2113), .in1(R8955), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2180 (.out1(_2080), .in1(R8957), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2163 (.out1(_2063), .in1(R8959), .in2(_2062));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2144 (.out1(_2044), .in1(R8960), .in2(63 'd 6148914691236517205));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2127 (.out1(_2027), .in1(R8962), .in2(1 'd 1));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op2094 (.out1(_1997), .in1(R8964), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2059 (.out1(_1962), .in1(_1944), .in2(_1961));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op2005 (.out1(_1911), .in1(R8967), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1970 (.out1(_1876), .in1(_1858), .in2(_1875));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op1916 (.out1(_1825), .in1(R8970), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1881 (.out1(_1790), .in1(_1772), .in2(_1789));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op1827 (.out1(_1739), .in1(R8973), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1792 (.out1(_1704), .in1(_1686), .in2(_1703));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op1738 (.out1(_1653), .in1(R8976), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1703 (.out1(_1618), .in1(_1600), .in2(_1617));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op1649 (.out1(_1567), .in1(R8979), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1614 (.out1(_1532), .in1(_1514), .in2(_1531));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op1560 (.out1(_1481), .in1(R8982), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1525 (.out1(_1446), .in1(_1428), .in2(_1445));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op1471 (.out1(_1395), .in1(R8985), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1436 (.out1(_1360), .in1(_1342), .in2(_1359));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op1382 (.out1(_1309), .in1(R8988), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1347 (.out1(_1274), .in1(_1256), .in2(_1273));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2590 (.out1(_2475), .in1(R8926), .in2(_2474));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2565 (.out1(_2450), .in1(R8907), .in2(R8928));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2501 (.out1(_2389), .in1(R8933), .in2(_2388));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2476 (.out1(_2364), .in1(R8908), .in2(R8935));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2412 (.out1(_2303), .in1(R8940), .in2(_2302));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2387 (.out1(_2278), .in1(R8909), .in2(R8942));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2323 (.out1(_2217), .in1(R8947), .in2(_2216));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2298 (.out1(_2192), .in1(R8910), .in2(R8949));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2234 (.out1(_2131), .in1(R8954), .in2(_2130));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2209 (.out1(_2106), .in1(R8911), .in2(R8956));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2145 (.out1(_2045), .in1(R8961), .in2(_2044));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2120 (.out1(_2020), .in1(R8912), .in2(R8963));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2557 (.out1(_2442), .in1(_2441), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2468 (.out1(_2356), .in1(_2355), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2379 (.out1(_2270), .in1(_2269), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2290 (.out1(_2184), .in1(_2183), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2201 (.out1(_2098), .in1(_2097), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2112 (.out1(_2012), .in1(_2011), .in2(2 'd 2));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2024 (.out1(_1927), .in1(b64_popcnt_2590_D), .in2(R8913));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1935 (.out1(_1841), .in1(b72_popcnt_2601_D), .in2(R8914));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1846 (.out1(_1755), .in1(b80_popcnt_2611_D), .in2(R8915));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1757 (.out1(_1669), .in1(b88_popcnt_2621_D), .in2(R8916));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1668 (.out1(_1583), .in1(b96_popcnt_2631_D), .in2(R8917));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1579 (.out1(_1497), .in1(b104_popcnt_2641_D), .in2(R8918));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1490 (.out1(_1411), .in1(b112_popcnt_2651_D), .in2(R8919));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1401 (.out1(_1325), .in1(b120_popcnt_2661_D), .in2(R8920));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1312 (.out1(_1239), .in1(b128_popcnt_2670_D), .in2(R8921));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2626 (.out1(_2511), .in1(_2510), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2609 (.out1(_2494), .in1(_2493), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2573 (.out1(_2458), .in1(_2457), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2537 (.out1(_2425), .in1(_2424), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2520 (.out1(_2408), .in1(_2407), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2484 (.out1(_2372), .in1(_2371), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2448 (.out1(_2339), .in1(_2338), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2431 (.out1(_2322), .in1(_2321), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2395 (.out1(_2286), .in1(_2285), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2359 (.out1(_2253), .in1(_2252), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2342 (.out1(_2236), .in1(_2235), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2306 (.out1(_2200), .in1(_2199), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2270 (.out1(_2167), .in1(_2166), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2253 (.out1(_2150), .in1(_2149), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2217 (.out1(_2114), .in1(_2113), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2181 (.out1(_2081), .in1(_2080), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2164 (.out1(_2064), .in1(_2063), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2128 (.out1(_2028), .in1(_2027), .in2(63 'd 6148914691236517205));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2095 (.out1(_1998), .in1(_1962), .in2(_1997));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2006 (.out1(_1912), .in1(_1876), .in2(_1911));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1917 (.out1(_1826), .in1(_1790), .in2(_1825));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1828 (.out1(_1740), .in1(_1704), .in2(_1739));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1739 (.out1(_1654), .in1(_1618), .in2(_1653));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1650 (.out1(_1568), .in1(_1532), .in2(_1567));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1561 (.out1(_1482), .in1(_1446), .in2(_1481));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1472 (.out1(_1396), .in1(_1360), .in2(_1395));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1383 (.out1(_1310), .in1(_1274), .in2(_1309));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2627 (.out1(_2512), .in1(_2494), .in2(_2511));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2591 (.out1(_2476), .in1(_2475), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2574 (.out1(_2459), .in1(_2450), .in2(_2458));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2538 (.out1(_2426), .in1(_2408), .in2(_2425));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2502 (.out1(_2390), .in1(_2389), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2485 (.out1(_2373), .in1(_2364), .in2(_2372));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2449 (.out1(_2340), .in1(_2322), .in2(_2339));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2413 (.out1(_2304), .in1(_2303), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2396 (.out1(_2287), .in1(_2278), .in2(_2286));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2360 (.out1(_2254), .in1(_2236), .in2(_2253));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2324 (.out1(_2218), .in1(_2217), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2307 (.out1(_2201), .in1(_2192), .in2(_2200));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2271 (.out1(_2168), .in1(_2150), .in2(_2167));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2235 (.out1(_2132), .in1(_2131), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2218 (.out1(_2115), .in1(_2106), .in2(_2114));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2182 (.out1(_2082), .in1(_2064), .in2(_2081));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2146 (.out1(_2046), .in1(_2045), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2129 (.out1(_2029), .in1(_2020), .in2(_2028));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op2096 (.out1(_1999), .in1(_1998), .in2(60 'd 1085102592571150095));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op2007 (.out1(_1913), .in1(_1912), .in2(60 'd 1085102592571150095));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op1918 (.out1(_1827), .in1(_1826), .in2(60 'd 1085102592571150095));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op1829 (.out1(_1741), .in1(_1740), .in2(60 'd 1085102592571150095));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op1740 (.out1(_1655), .in1(_1654), .in2(60 'd 1085102592571150095));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op1651 (.out1(_1569), .in1(_1568), .in2(60 'd 1085102592571150095));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op1562 (.out1(_1483), .in1(_1482), .in2(60 'd 1085102592571150095));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op1473 (.out1(_1397), .in1(_1396), .in2(60 'd 1085102592571150095));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op1384 (.out1(_1311), .in1(_1310), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3285 (.out1(R3286), .clock(clock), .in1(R3285));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3912 (.out1(R3913), .clock(clock), .in1(R3912));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4497 (.out1(R4498), .clock(clock), .in1(R4497));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5040 (.out1(R5041), .clock(clock), .in1(R5040));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5541 (.out1(R5542), .clock(clock), .in1(R5541));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6000 (.out1(R6001), .clock(clock), .in1(R6000));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6414 (.out1(R6415), .clock(clock), .in1(R6414));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6787 (.out1(R6788), .clock(clock), .in1(R6787));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7117 (.out1(R7118), .clock(clock), .in1(R7117));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7405 (.out1(R7406), .clock(clock), .in1(R7405));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7651 (.out1(R7652), .clock(clock), .in1(R7651));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7855 (.out1(R7856), .clock(clock), .in1(R7855));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8017 (.out1(R8018), .clock(clock), .in1(R8017));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8137 (.out1(R8138), .clock(clock), .in1(R8137));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8264 (.out1(R8265), .clock(clock), .in1(R8264));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8275 (.out1(R8276), .clock(clock), .in1(R8275));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8286 (.out1(R8287), .clock(clock), .in1(R8286));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8297 (.out1(R8298), .clock(clock), .in1(R8297));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8308 (.out1(R8309), .clock(clock), .in1(R8308));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8319 (.out1(R8320), .clock(clock), .in1(R8319));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8330 (.out1(R8331), .clock(clock), .in1(R8330));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8341 (.out1(R8342), .clock(clock), .in1(R8341));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8352 (.out1(R8353), .clock(clock), .in1(R8352));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8377 (.out1(R8378), .clock(clock), .in1(R8377));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8388 (.out1(R8389), .clock(clock), .in1(R8388));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8399 (.out1(R8400), .clock(clock), .in1(R8399));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8410 (.out1(R8411), .clock(clock), .in1(R8410));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8421 (.out1(R8422), .clock(clock), .in1(R8421));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8432 (.out1(R8433), .clock(clock), .in1(R8432));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8990 (.out1(R8991), .clock(clock), .in1(_2442));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8991 (.out1(R8992), .clock(clock), .in1(_2356));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8992 (.out1(R8993), .clock(clock), .in1(_2270));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8993 (.out1(R8994), .clock(clock), .in1(_2184));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8994 (.out1(R8995), .clock(clock), .in1(_2098));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8995 (.out1(R8996), .clock(clock), .in1(_2012));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8996 (.out1(R8997), .clock(clock), .in1(_1927));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8997 (.out1(R8998), .clock(clock), .in1(_1841));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8998 (.out1(R8999), .clock(clock), .in1(_1755));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8999 (.out1(R9000), .clock(clock), .in1(_1669));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9000 (.out1(R9001), .clock(clock), .in1(_1583));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9001 (.out1(R9002), .clock(clock), .in1(_1497));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9002 (.out1(R9003), .clock(clock), .in1(_1411));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9003 (.out1(R9004), .clock(clock), .in1(_1325));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9004 (.out1(R9005), .clock(clock), .in1(_1239));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9005 (.out1(R9006), .clock(clock), .in1(_2512));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9006 (.out1(R9007), .clock(clock), .in1(_2476));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9007 (.out1(R9008), .clock(clock), .in1(_2459));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9008 (.out1(R9009), .clock(clock), .in1(_2426));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9009 (.out1(R9010), .clock(clock), .in1(_2390));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9010 (.out1(R9011), .clock(clock), .in1(_2373));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9011 (.out1(R9012), .clock(clock), .in1(_2340));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9012 (.out1(R9013), .clock(clock), .in1(_2304));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9013 (.out1(R9014), .clock(clock), .in1(_2287));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9014 (.out1(R9015), .clock(clock), .in1(_2254));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9015 (.out1(R9016), .clock(clock), .in1(_2218));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9016 (.out1(R9017), .clock(clock), .in1(_2201));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9017 (.out1(R9018), .clock(clock), .in1(_2168));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9018 (.out1(R9019), .clock(clock), .in1(_2132));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9019 (.out1(R9020), .clock(clock), .in1(_2115));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9020 (.out1(R9021), .clock(clock), .in1(_2082));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9021 (.out1(R9022), .clock(clock), .in1(_2046));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9022 (.out1(R9023), .clock(clock), .in1(_2029));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9023 (.out1(R9024), .clock(clock), .in1(_1999));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9024 (.out1(R9025), .clock(clock), .in1(_1913));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9025 (.out1(R9026), .clock(clock), .in1(_1827));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9026 (.out1(R9027), .clock(clock), .in1(_1741));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9027 (.out1(R9028), .clock(clock), .in1(_1655));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9028 (.out1(R9029), .clock(clock), .in1(_1569));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9029 (.out1(R9030), .clock(clock), .in1(_1483));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9030 (.out1(R9031), .clock(clock), .in1(_1397));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9031 (.out1(R9032), .clock(clock), .in1(_1311));
  SRAM op2025 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1928),.ADR(R8997));
  SRAM op1936 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1842),.ADR(R8998));
  SRAM op1847 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1756),.ADR(R8999));
  SRAM op1758 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1670),.ADR(R9000));
  SRAM op1669 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1584),.ADR(R9001));
  SRAM op1580 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1498),.ADR(R9002));
  SRAM op1491 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1412),.ADR(R9003));
  SRAM op1402 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1326),.ADR(R9004));
  SRAM op1313 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1240),.ADR(R9005));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op2097 (.out1(_2000), .in1(R9024), .in2(57 'd 72340172838076673));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op2008 (.out1(_1914), .in1(R9025), .in2(57 'd 72340172838076673));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op1919 (.out1(_1828), .in1(R9026), .in2(57 'd 72340172838076673));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op1830 (.out1(_1742), .in1(R9027), .in2(57 'd 72340172838076673));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op1741 (.out1(_1656), .in1(R9028), .in2(57 'd 72340172838076673));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op1652 (.out1(_1570), .in1(R9029), .in2(57 'd 72340172838076673));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op1563 (.out1(_1484), .in1(R9030), .in2(57 'd 72340172838076673));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op1474 (.out1(_1398), .in1(R9031), .in2(57 'd 72340172838076673));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op1385 (.out1(_1312), .in1(R9032), .in2(57 'd 72340172838076673));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2592 (.out1(_2477), .in1(R9007), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2575 (.out1(_2460), .in1(R9008), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2503 (.out1(_2391), .in1(R9010), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2486 (.out1(_2374), .in1(R9011), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2414 (.out1(_2305), .in1(R9013), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2397 (.out1(_2288), .in1(R9014), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2325 (.out1(_2219), .in1(R9016), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2308 (.out1(_2202), .in1(R9017), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2236 (.out1(_2133), .in1(R9019), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2219 (.out1(_2116), .in1(R9020), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2147 (.out1(_2047), .in1(R9022), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2130 (.out1(_2030), .in1(R9023), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op2628 (.out1(_2513), .in1(R9006), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2593 (.out1(_2478), .in1(_2460), .in2(_2477));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op2539 (.out1(_2427), .in1(R9009), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2504 (.out1(_2392), .in1(_2374), .in2(_2391));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op2450 (.out1(_2341), .in1(R9012), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2415 (.out1(_2306), .in1(_2288), .in2(_2305));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op2361 (.out1(_2255), .in1(R9015), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2326 (.out1(_2220), .in1(_2202), .in2(_2219));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op2272 (.out1(_2169), .in1(R9018), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2237 (.out1(_2134), .in1(_2116), .in2(_2133));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op2183 (.out1(_2083), .in1(R9021), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2148 (.out1(_2048), .in1(_2030), .in2(_2047));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2558 (.out1(_2443), .in1(b16_popcnt_2529_D), .in2(R8991));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2469 (.out1(_2357), .in1(b24_popcnt_2540_D), .in2(R8992));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2380 (.out1(_2271), .in1(b32_popcnt_2550_D), .in2(R8993));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2291 (.out1(_2185), .in1(b40_popcnt_2560_D), .in2(R8994));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2202 (.out1(_2099), .in1(b48_popcnt_2570_D), .in2(R8995));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2113 (.out1(_2013), .in1(b56_popcnt_2580_D), .in2(R8996));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2629 (.out1(_2514), .in1(_2478), .in2(_2513));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2540 (.out1(_2428), .in1(_2392), .in2(_2427));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2451 (.out1(_2342), .in1(_2306), .in2(_2341));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2362 (.out1(_2256), .in1(_2220), .in2(_2255));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2273 (.out1(_2170), .in1(_2134), .in2(_2169));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2184 (.out1(_2084), .in1(_2048), .in2(_2083));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op2630 (.out1(_2515), .in1(_2514), .in2(60 'd 1085102592571150095));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op2541 (.out1(_2429), .in1(_2428), .in2(60 'd 1085102592571150095));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op2452 (.out1(_2343), .in1(_2342), .in2(60 'd 1085102592571150095));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op2363 (.out1(_2257), .in1(_2256), .in2(60 'd 1085102592571150095));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op2274 (.out1(_2171), .in1(_2170), .in2(60 'd 1085102592571150095));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op2185 (.out1(_2085), .in1(_2084), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3286 (.out1(R3287), .clock(clock), .in1(R3286));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3913 (.out1(R3914), .clock(clock), .in1(R3913));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4498 (.out1(R4499), .clock(clock), .in1(R4498));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5041 (.out1(R5042), .clock(clock), .in1(R5041));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5542 (.out1(R5543), .clock(clock), .in1(R5542));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6001 (.out1(R6002), .clock(clock), .in1(R6001));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6415 (.out1(R6416), .clock(clock), .in1(R6415));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6788 (.out1(R6789), .clock(clock), .in1(R6788));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7118 (.out1(R7119), .clock(clock), .in1(R7118));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7406 (.out1(R7407), .clock(clock), .in1(R7406));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7652 (.out1(R7653), .clock(clock), .in1(R7652));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7856 (.out1(R7857), .clock(clock), .in1(R7856));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8018 (.out1(R8019), .clock(clock), .in1(R8018));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8138 (.out1(R8139), .clock(clock), .in1(R8138));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8265 (.out1(R8266), .clock(clock), .in1(R8265));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8276 (.out1(R8277), .clock(clock), .in1(R8276));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8287 (.out1(R8288), .clock(clock), .in1(R8287));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8298 (.out1(R8299), .clock(clock), .in1(R8298));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8309 (.out1(R8310), .clock(clock), .in1(R8309));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8320 (.out1(R8321), .clock(clock), .in1(R8320));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8331 (.out1(R8332), .clock(clock), .in1(R8331));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8342 (.out1(R8343), .clock(clock), .in1(R8342));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8353 (.out1(R8354), .clock(clock), .in1(R8353));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8378 (.out1(R8379), .clock(clock), .in1(R8378));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8389 (.out1(R8390), .clock(clock), .in1(R8389));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8400 (.out1(R8401), .clock(clock), .in1(R8400));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8411 (.out1(R8412), .clock(clock), .in1(R8411));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8422 (.out1(R8423), .clock(clock), .in1(R8422));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8433 (.out1(R8434), .clock(clock), .in1(R8433));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9032 (.out1(R9033), .clock(clock), .in1(_1928));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9033 (.out1(R9034), .clock(clock), .in1(_1842));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9034 (.out1(R9035), .clock(clock), .in1(_1756));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9035 (.out1(R9036), .clock(clock), .in1(_1670));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9036 (.out1(R9037), .clock(clock), .in1(_1584));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9037 (.out1(R9038), .clock(clock), .in1(_1498));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9038 (.out1(R9039), .clock(clock), .in1(_1412));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9039 (.out1(R9040), .clock(clock), .in1(_1326));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9040 (.out1(R9041), .clock(clock), .in1(_1240));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9041 (.out1(R9042), .clock(clock), .in1(_2000));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9042 (.out1(R9043), .clock(clock), .in1(_1914));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9043 (.out1(R9044), .clock(clock), .in1(_1828));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9044 (.out1(R9045), .clock(clock), .in1(_1742));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9045 (.out1(R9046), .clock(clock), .in1(_1656));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9046 (.out1(R9047), .clock(clock), .in1(_1570));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9047 (.out1(R9048), .clock(clock), .in1(_1484));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9048 (.out1(R9049), .clock(clock), .in1(_1398));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9049 (.out1(R9050), .clock(clock), .in1(_1312));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9050 (.out1(R9051), .clock(clock), .in1(_2443));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9051 (.out1(R9052), .clock(clock), .in1(_2357));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9052 (.out1(R9053), .clock(clock), .in1(_2271));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9053 (.out1(R9054), .clock(clock), .in1(_2185));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9054 (.out1(R9055), .clock(clock), .in1(_2099));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9055 (.out1(R9056), .clock(clock), .in1(_2013));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9056 (.out1(R9057), .clock(clock), .in1(_2515));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9057 (.out1(R9058), .clock(clock), .in1(_2429));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9058 (.out1(R9059), .clock(clock), .in1(_2343));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9059 (.out1(R9060), .clock(clock), .in1(_2257));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9060 (.out1(R9061), .clock(clock), .in1(_2171));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9061 (.out1(R9062), .clock(clock), .in1(_2085));
  SRAM op2559 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2444),.ADR(R9051));
  SRAM op2470 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2358),.ADR(R9052));
  SRAM op2381 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2272),.ADR(R9053));
  SRAM op2292 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2186),.ADR(R9054));
  SRAM op2203 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2100),.ADR(R9055));
  SRAM op2114 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2014),.ADR(R9056));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op2631 (.out1(_2516), .in1(R9057), .in2(57 'd 72340172838076673));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op2542 (.out1(_2430), .in1(R9058), .in2(57 'd 72340172838076673));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op2453 (.out1(_2344), .in1(R9059), .in2(57 'd 72340172838076673));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op2364 (.out1(_2258), .in1(R9060), .in2(57 'd 72340172838076673));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op2275 (.out1(_2172), .in1(R9061), .in2(57 'd 72340172838076673));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op2186 (.out1(_2086), .in1(R9062), .in2(57 'd 72340172838076673));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op2098 (.out1(_2001), .in1(R9042), .in2(6 'd 56));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op2009 (.out1(_1915), .in1(R9043), .in2(6 'd 56));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op1920 (.out1(_1829), .in1(R9044), .in2(6 'd 56));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op1831 (.out1(_1743), .in1(R9045), .in2(6 'd 56));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op1742 (.out1(_1657), .in1(R9046), .in2(6 'd 56));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op1653 (.out1(_1571), .in1(R9047), .in2(6 'd 56));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op1564 (.out1(_1485), .in1(R9048), .in2(6 'd 56));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op1475 (.out1(_1399), .in1(R9049), .in2(6 'd 56));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op1386 (.out1(_1313), .in1(R9050), .in2(6 'd 56));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op2099 (.out1(_2002), .in1(_2001));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op2010 (.out1(_1916), .in1(_1915));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1921 (.out1(_1830), .in1(_1829));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1832 (.out1(_1744), .in1(_1743));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1743 (.out1(_1658), .in1(_1657));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1654 (.out1(_1572), .in1(_1571));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1565 (.out1(_1486), .in1(_1485));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1476 (.out1(_1400), .in1(_1399));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1387 (.out1(_1314), .in1(_1313));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2100 (.out1(n_idx_2591), .in1(R9033), .in2(_2002));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2011 (.out1(n_idx_2602), .in1(R9034), .in2(_1916));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1922 (.out1(n_idx_2612), .in1(R9035), .in2(_1830));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1833 (.out1(n_idx_2622), .in1(R9036), .in2(_1744));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1744 (.out1(n_idx_2632), .in1(R9037), .in2(_1658));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1655 (.out1(n_idx_2642), .in1(R9038), .in2(_1572));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1566 (.out1(n_idx_2652), .in1(R9039), .in2(_1486));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1477 (.out1(n_idx_2662), .in1(R9040), .in2(_1400));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1388 (.out1(n_idx_2671), .in1(R9041), .in2(_1314));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3287 (.out1(R3288), .clock(clock), .in1(R3287));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3914 (.out1(R3915), .clock(clock), .in1(R3914));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4499 (.out1(R4500), .clock(clock), .in1(R4499));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5042 (.out1(R5043), .clock(clock), .in1(R5042));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5543 (.out1(R5544), .clock(clock), .in1(R5543));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6002 (.out1(R6003), .clock(clock), .in1(R6002));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6416 (.out1(R6417), .clock(clock), .in1(R6416));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6789 (.out1(R6790), .clock(clock), .in1(R6789));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7119 (.out1(R7120), .clock(clock), .in1(R7119));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7407 (.out1(R7408), .clock(clock), .in1(R7407));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7653 (.out1(R7654), .clock(clock), .in1(R7653));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7857 (.out1(R7858), .clock(clock), .in1(R7857));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8019 (.out1(R8020), .clock(clock), .in1(R8019));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8139 (.out1(R8140), .clock(clock), .in1(R8139));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8266 (.out1(R8267), .clock(clock), .in1(R8266));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8277 (.out1(R8278), .clock(clock), .in1(R8277));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8288 (.out1(R8289), .clock(clock), .in1(R8288));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8299 (.out1(R8300), .clock(clock), .in1(R8299));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8310 (.out1(R8311), .clock(clock), .in1(R8310));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8321 (.out1(R8322), .clock(clock), .in1(R8321));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8332 (.out1(R8333), .clock(clock), .in1(R8332));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8343 (.out1(R8344), .clock(clock), .in1(R8343));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8354 (.out1(R8355), .clock(clock), .in1(R8354));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8379 (.out1(R8380), .clock(clock), .in1(R8379));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8390 (.out1(R8391), .clock(clock), .in1(R8390));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8401 (.out1(R8402), .clock(clock), .in1(R8401));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8412 (.out1(R8413), .clock(clock), .in1(R8412));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8423 (.out1(R8424), .clock(clock), .in1(R8423));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8434 (.out1(R8435), .clock(clock), .in1(R8434));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9062 (.out1(R9063), .clock(clock), .in1(_2444));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9063 (.out1(R9064), .clock(clock), .in1(_2358));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9064 (.out1(R9065), .clock(clock), .in1(_2272));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9065 (.out1(R9066), .clock(clock), .in1(_2186));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9066 (.out1(R9067), .clock(clock), .in1(_2100));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9067 (.out1(R9068), .clock(clock), .in1(_2014));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9068 (.out1(R9069), .clock(clock), .in1(_2516));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9069 (.out1(R9070), .clock(clock), .in1(_2430));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9070 (.out1(R9071), .clock(clock), .in1(_2344));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9071 (.out1(R9072), .clock(clock), .in1(_2258));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9072 (.out1(R9073), .clock(clock), .in1(_2172));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9073 (.out1(R9074), .clock(clock), .in1(_2086));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9074 (.out1(R9075), .clock(clock), .in1(n_idx_2591));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9075 (.out1(R9076), .clock(clock), .in1(n_idx_2602));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9076 (.out1(R9077), .clock(clock), .in1(n_idx_2612));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9077 (.out1(R9078), .clock(clock), .in1(n_idx_2622));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9078 (.out1(R9079), .clock(clock), .in1(n_idx_2632));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9079 (.out1(R9080), .clock(clock), .in1(n_idx_2642));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9080 (.out1(R9081), .clock(clock), .in1(n_idx_2652));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9081 (.out1(R9082), .clock(clock), .in1(n_idx_2662));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9082 (.out1(R9083), .clock(clock), .in1(n_idx_2671));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op2632 (.out1(_2517), .in1(R9069), .in2(6 'd 56));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op2543 (.out1(_2431), .in1(R9070), .in2(6 'd 56));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op2454 (.out1(_2345), .in1(R9071), .in2(6 'd 56));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op2365 (.out1(_2259), .in1(R9072), .in2(6 'd 56));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op2276 (.out1(_2173), .in1(R9073), .in2(6 'd 56));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op2187 (.out1(_2087), .in1(R9074), .in2(6 'd 56));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2101 (.out1(_2003), .in1(R9075));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2012 (.out1(_1917), .in1(R9076));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1923 (.out1(_1831), .in1(R9077));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1834 (.out1(_1745), .in1(R9078));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1745 (.out1(_1659), .in1(R9079));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1656 (.out1(_1573), .in1(R9080));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1567 (.out1(_1487), .in1(R9081));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1478 (.out1(_1401), .in1(R9082));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1389 (.out1(_1315), .in1(R9083));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2102 (.out1(_2004), .in1(leafN_2531_D), .in2(_2003));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2013 (.out1(_1918), .in1(leafN_2531_D), .in2(_1917));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1924 (.out1(_1832), .in1(leafN_2531_D), .in2(_1831));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1835 (.out1(_1746), .in1(leafN_2531_D), .in2(_1745));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1746 (.out1(_1660), .in1(leafN_2531_D), .in2(_1659));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1657 (.out1(_1574), .in1(leafN_2531_D), .in2(_1573));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1568 (.out1(_1488), .in1(leafN_2531_D), .in2(_1487));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1479 (.out1(_1402), .in1(leafN_2531_D), .in2(_1401));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1390 (.out1(_1316), .in1(leafN_2531_D), .in2(_1315));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op2633 (.out1(_2518), .in1(_2517));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op2544 (.out1(_2432), .in1(_2431));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op2455 (.out1(_2346), .in1(_2345));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op2366 (.out1(_2260), .in1(_2259));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op2277 (.out1(_2174), .in1(_2173));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op2188 (.out1(_2088), .in1(_2087));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2634 (.out1(n_idx_2530), .in1(R9063), .in2(_2518));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2545 (.out1(n_idx_2541), .in1(R9064), .in2(_2432));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2456 (.out1(n_idx_2551), .in1(R9065), .in2(_2346));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2367 (.out1(n_idx_2561), .in1(R9066), .in2(_2260));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2278 (.out1(n_idx_2571), .in1(R9067), .in2(_2174));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2189 (.out1(n_idx_2581), .in1(R9068), .in2(_2088));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3288 (.out1(R3289), .clock(clock), .in1(R3288));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3915 (.out1(R3916), .clock(clock), .in1(R3915));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4500 (.out1(R4501), .clock(clock), .in1(R4500));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5043 (.out1(R5044), .clock(clock), .in1(R5043));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5544 (.out1(R5545), .clock(clock), .in1(R5544));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6003 (.out1(R6004), .clock(clock), .in1(R6003));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6417 (.out1(R6418), .clock(clock), .in1(R6417));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6790 (.out1(R6791), .clock(clock), .in1(R6790));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7120 (.out1(R7121), .clock(clock), .in1(R7120));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7408 (.out1(R7409), .clock(clock), .in1(R7408));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7654 (.out1(R7655), .clock(clock), .in1(R7654));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7858 (.out1(R7859), .clock(clock), .in1(R7858));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8020 (.out1(R8021), .clock(clock), .in1(R8020));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8140 (.out1(R8141), .clock(clock), .in1(R8140));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8267 (.out1(R8268), .clock(clock), .in1(R8267));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8278 (.out1(R8279), .clock(clock), .in1(R8278));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8289 (.out1(R8290), .clock(clock), .in1(R8289));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8300 (.out1(R8301), .clock(clock), .in1(R8300));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8311 (.out1(R8312), .clock(clock), .in1(R8311));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8322 (.out1(R8323), .clock(clock), .in1(R8322));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8333 (.out1(R8334), .clock(clock), .in1(R8333));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8344 (.out1(R8345), .clock(clock), .in1(R8344));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8355 (.out1(R8356), .clock(clock), .in1(R8355));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8380 (.out1(R8381), .clock(clock), .in1(R8380));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8391 (.out1(R8392), .clock(clock), .in1(R8391));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8402 (.out1(R8403), .clock(clock), .in1(R8402));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8413 (.out1(R8414), .clock(clock), .in1(R8413));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8424 (.out1(R8425), .clock(clock), .in1(R8424));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8435 (.out1(R8436), .clock(clock), .in1(R8435));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9083 (.out1(R9084), .clock(clock), .in1(_2004));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9084 (.out1(R9085), .clock(clock), .in1(_1918));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9085 (.out1(R9086), .clock(clock), .in1(_1832));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9086 (.out1(R9087), .clock(clock), .in1(_1746));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9087 (.out1(R9088), .clock(clock), .in1(_1660));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9088 (.out1(R9089), .clock(clock), .in1(_1574));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9089 (.out1(R9090), .clock(clock), .in1(_1488));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9090 (.out1(R9091), .clock(clock), .in1(_1402));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9091 (.out1(R9092), .clock(clock), .in1(_1316));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9092 (.out1(R9093), .clock(clock), .in1(n_idx_2530));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9093 (.out1(R9094), .clock(clock), .in1(n_idx_2541));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9094 (.out1(R9095), .clock(clock), .in1(n_idx_2551));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9095 (.out1(R9096), .clock(clock), .in1(n_idx_2561));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9096 (.out1(R9097), .clock(clock), .in1(n_idx_2571));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9097 (.out1(R9098), .clock(clock), .in1(n_idx_2581));
  SRAM op2103 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2592),.ADR(R9084));
  SRAM op2014 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2603),.ADR(R9085));
  SRAM op1925 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2613),.ADR(R9086));
  SRAM op1836 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2623),.ADR(R9087));
  SRAM op1747 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2633),.ADR(R9088));
  SRAM op1658 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2643),.ADR(R9089));
  SRAM op1569 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2653),.ADR(R9090));
  SRAM op1480 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2663),.ADR(R9091));
  SRAM op1391 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2672),.ADR(R9092));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2635 (.out1(_2519), .in1(R9093));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2546 (.out1(_2433), .in1(R9094));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2457 (.out1(_2347), .in1(R9095));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2368 (.out1(_2261), .in1(R9096));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2279 (.out1(_2175), .in1(R9097));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2190 (.out1(_2089), .in1(R9098));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2636 (.out1(_2520), .in1(leafN_2531_D), .in2(_2519));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2547 (.out1(_2434), .in1(leafN_2531_D), .in2(_2433));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2458 (.out1(_2348), .in1(leafN_2531_D), .in2(_2347));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2369 (.out1(_2262), .in1(leafN_2531_D), .in2(_2261));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2280 (.out1(_2176), .in1(leafN_2531_D), .in2(_2175));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2191 (.out1(_2090), .in1(leafN_2531_D), .in2(_2089));
  cast #(.BITSIZE_in1(1), .BITSIZE_out1(8)) op2638 (.out1(_2673), .in1(1 'd 1));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3289 (.out1(R3290), .clock(clock), .in1(R3289));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3916 (.out1(R3917), .clock(clock), .in1(R3916));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4501 (.out1(R4502), .clock(clock), .in1(R4501));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5044 (.out1(R5045), .clock(clock), .in1(R5044));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5545 (.out1(R5546), .clock(clock), .in1(R5545));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6004 (.out1(R6005), .clock(clock), .in1(R6004));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6418 (.out1(R6419), .clock(clock), .in1(R6418));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6791 (.out1(R6792), .clock(clock), .in1(R6791));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7121 (.out1(R7122), .clock(clock), .in1(R7121));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7409 (.out1(R7410), .clock(clock), .in1(R7409));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7655 (.out1(R7656), .clock(clock), .in1(R7655));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7859 (.out1(R7860), .clock(clock), .in1(R7859));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8021 (.out1(R8022), .clock(clock), .in1(R8021));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8141 (.out1(R8142), .clock(clock), .in1(R8141));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8268 (.out1(R8269), .clock(clock), .in1(R8268));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8279 (.out1(R8280), .clock(clock), .in1(R8279));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8290 (.out1(R8291), .clock(clock), .in1(R8290));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8301 (.out1(R8302), .clock(clock), .in1(R8301));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8312 (.out1(R8313), .clock(clock), .in1(R8312));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8323 (.out1(R8324), .clock(clock), .in1(R8323));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8334 (.out1(R8335), .clock(clock), .in1(R8334));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8345 (.out1(R8346), .clock(clock), .in1(R8345));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8356 (.out1(R8357), .clock(clock), .in1(R8356));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8381 (.out1(R8382), .clock(clock), .in1(R8381));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8392 (.out1(R8393), .clock(clock), .in1(R8392));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8403 (.out1(R8404), .clock(clock), .in1(R8403));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8414 (.out1(R8415), .clock(clock), .in1(R8414));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8425 (.out1(R8426), .clock(clock), .in1(R8425));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8436 (.out1(R8437), .clock(clock), .in1(R8436));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op9098 (.out1(R9099), .clock(clock), .in1(_2592));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op9099 (.out1(R9100), .clock(clock), .in1(_2603));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op9100 (.out1(R9101), .clock(clock), .in1(_2613));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op9101 (.out1(R9102), .clock(clock), .in1(_2623));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op9102 (.out1(R9103), .clock(clock), .in1(_2633));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op9103 (.out1(R9104), .clock(clock), .in1(_2643));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op9104 (.out1(R9105), .clock(clock), .in1(_2653));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op9105 (.out1(R9106), .clock(clock), .in1(_2663));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op9106 (.out1(R9107), .clock(clock), .in1(_2672));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9107 (.out1(R9108), .clock(clock), .in1(_2520));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9108 (.out1(R9109), .clock(clock), .in1(_2434));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9109 (.out1(R9110), .clock(clock), .in1(_2348));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9110 (.out1(R9111), .clock(clock), .in1(_2262));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9111 (.out1(R9112), .clock(clock), .in1(_2176));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9112 (.out1(R9113), .clock(clock), .in1(_2090));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op9113 (.out1(R9114), .clock(clock), .in1(_2673));
  SRAM op2637 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2532),.ADR(R9108));
  SRAM op2548 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2542),.ADR(R9109));
  SRAM op2459 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2552),.ADR(R9110));
  SRAM op2370 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2562),.ADR(R9111));
  SRAM op2281 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2572),.ADR(R9112));
  SRAM op2192 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2582),.ADR(R9113));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op2652 (.out1(mux13), .in1(R9114), .in2(R9106), .sel(R8346));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op2653 (.out1(mux14), .in1(R9114), .in2(R9107), .sel(R8357));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op2651 (.out1(mux12), .in1(R9114), .in2(R9105), .sel(R8335));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op2654 (.out1(mux15), .in1(mux13), .in2(mux14), .sel(R8142));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op2650 (.out1(mux11), .in1(R9114), .in2(R9104), .sel(R8324));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op2655 (.out1(mux16), .in1(mux12), .in2(mux15), .sel(R8022));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op2649 (.out1(mux10), .in1(R9114), .in2(R9103), .sel(R8313));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op2656 (.out1(mux17), .in1(mux11), .in2(mux16), .sel(R7860));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op2648 (.out1(mux9), .in1(R9114), .in2(R9102), .sel(R8302));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op2657 (.out1(mux18), .in1(mux10), .in2(mux17), .sel(R7656));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op2647 (.out1(mux8), .in1(R9114), .in2(R9101), .sel(R8291));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op2658 (.out1(mux19), .in1(mux9), .in2(mux18), .sel(R7410));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op2646 (.out1(mux7), .in1(R9114), .in2(R9100), .sel(R8280));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op2659 (.out1(mux20), .in1(mux8), .in2(mux19), .sel(R7122));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op2645 (.out1(mux6), .in1(R9114), .in2(R9099), .sel(R8269));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op2660 (.out1(mux21), .in1(mux7), .in2(mux20), .sel(R6792));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3290 (.out1(R3291), .clock(clock), .in1(R3290));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3917 (.out1(R3918), .clock(clock), .in1(R3917));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4502 (.out1(R4503), .clock(clock), .in1(R4502));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5045 (.out1(R5046), .clock(clock), .in1(R5045));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5546 (.out1(R5547), .clock(clock), .in1(R5546));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6005 (.out1(R6006), .clock(clock), .in1(R6005));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6419 (.out1(R6420), .clock(clock), .in1(R6419));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8382 (.out1(R8383), .clock(clock), .in1(R8382));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8393 (.out1(R8394), .clock(clock), .in1(R8393));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8404 (.out1(R8405), .clock(clock), .in1(R8404));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8415 (.out1(R8416), .clock(clock), .in1(R8415));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8426 (.out1(R8427), .clock(clock), .in1(R8426));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8437 (.out1(R8438), .clock(clock), .in1(R8437));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op9114 (.out1(R9115), .clock(clock), .in1(R9114));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op9115 (.out1(R9116), .clock(clock), .in1(_2532));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op9116 (.out1(R9117), .clock(clock), .in1(_2542));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op9117 (.out1(R9118), .clock(clock), .in1(_2552));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op9118 (.out1(R9119), .clock(clock), .in1(_2562));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op9119 (.out1(R9120), .clock(clock), .in1(_2572));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op9120 (.out1(R9121), .clock(clock), .in1(_2582));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op9121 (.out1(R9122), .clock(clock), .in1(mux6));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op9122 (.out1(R9123), .clock(clock), .in1(mux21));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op2644 (.out1(mux5), .in1(R9115), .in2(R9121), .sel(R8438));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op2661 (.out1(mux22), .in1(R9122), .in2(R9123), .sel(R6420));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op2643 (.out1(mux4), .in1(R9115), .in2(R9120), .sel(R8427));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op2662 (.out1(mux23), .in1(mux5), .in2(mux22), .sel(R6006));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op2642 (.out1(mux3), .in1(R9115), .in2(R9119), .sel(R8416));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op2663 (.out1(mux24), .in1(mux4), .in2(mux23), .sel(R5547));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op2641 (.out1(mux2), .in1(R9115), .in2(R9118), .sel(R8405));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op2664 (.out1(mux25), .in1(mux3), .in2(mux24), .sel(R5046));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op2640 (.out1(mux1), .in1(R9115), .in2(R9117), .sel(R8394));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op2665 (.out1(mux26), .in1(mux2), .in2(mux25), .sel(R4503));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op2639 (.out1(mux0), .in1(R9115), .in2(R9116), .sel(R8383));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op2666 (.out1(mux27), .in1(mux1), .in2(mux26), .sel(R3918));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op2667 (.out1(mux28), .in1(mux0), .in2(mux27), .sel(R3291));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op9123 (.out1(R9124), .clock(clock), .in1(mux28));
endmodule