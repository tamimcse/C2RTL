`include "module_library.v"
`include "macros.v"

`timescale 1ns / 1ps
module top(clock, N16_3534_D, base1_16_3540_D, leafvec16_3539_D, base1_22_3549_D, leafvec22_3548_D, base1_28_3557_D, leafvec28_3556_D, base1_34_3565_D, leafvec34_3564_D, base1_40_3573_D, leafvec40_3572_D, base1_46_3581_D, leafvec46_3580_D, base1_52_3589_D, leafvec52_3588_D, base1_58_3597_D, leafvec58_3596_D, base1_64_3606_D, leafvec64_3605_D, base1_70_3614_D, leafvec70_3613_D, base1_76_3622_D, leafvec76_3621_D, base1_82_3630_D, leafvec82_3629_D, base1_88_3638_D, leafvec88_3637_D, base1_94_3646_D, leafvec94_3645_D, base1_100_3654_D, leafvec100_3653_D, base1_106_3662_D, leafvec106_3661_D, base1_112_3670_D, leafvec112_3669_D, base1_118_3678_D, leafvec118_3677_D, leafN_3542_D, base1_124_3685_D, leafvec124_3684_D, base0_118_3681_D, vec118_3676_D, base0_112_3673_D, vec112_3668_D, base0_106_3665_D, vec106_3660_D, base0_100_3657_D, vec100_3652_D, base0_94_3649_D, vec94_3644_D, base0_88_3641_D, vec88_3636_D, base0_82_3633_D, vec82_3628_D, base0_76_3625_D, vec76_3620_D, base0_70_3617_D, vec70_3612_D, base0_64_3609_D, vec64_3604_D, ip2_3602_D, base0_58_3600_D, vec58_3595_D, base0_52_3592_D, vec52_3587_D, base0_46_3584_D, vec46_3579_D, base0_40_3576_D, vec40_3571_D, base0_34_3568_D, vec34_3563_D, base0_28_3560_D, vec28_3555_D, base0_22_3552_D, vec22_3547_D, base0_16_3544_D, vec16_3538_D, dirC_3532_D, ip1_3530_D, R13573);
  //IN
  input clock;
  input [63:0] N16_3534_D;
  input [63:0] base1_16_3540_D;
  input [63:0] leafvec16_3539_D;
  input [63:0] base1_22_3549_D;
  input [63:0] leafvec22_3548_D;
  input [63:0] base1_28_3557_D;
  input [63:0] leafvec28_3556_D;
  input [63:0] base1_34_3565_D;
  input [63:0] leafvec34_3564_D;
  input [63:0] base1_40_3573_D;
  input [63:0] leafvec40_3572_D;
  input [63:0] base1_46_3581_D;
  input [63:0] leafvec46_3580_D;
  input [63:0] base1_52_3589_D;
  input [63:0] leafvec52_3588_D;
  input [63:0] base1_58_3597_D;
  input [63:0] leafvec58_3596_D;
  input [63:0] base1_64_3606_D;
  input [63:0] leafvec64_3605_D;
  input [63:0] base1_70_3614_D;
  input [63:0] leafvec70_3613_D;
  input [63:0] base1_76_3622_D;
  input [63:0] leafvec76_3621_D;
  input [63:0] base1_82_3630_D;
  input [63:0] leafvec82_3629_D;
  input [63:0] base1_88_3638_D;
  input [63:0] leafvec88_3637_D;
  input [63:0] base1_94_3646_D;
  input [63:0] leafvec94_3645_D;
  input [63:0] base1_100_3654_D;
  input [63:0] leafvec100_3653_D;
  input [63:0] base1_106_3662_D;
  input [63:0] leafvec106_3661_D;
  input [63:0] base1_112_3670_D;
  input [63:0] leafvec112_3669_D;
  input [63:0] base1_118_3678_D;
  input [63:0] leafvec118_3677_D;
  input [63:0] leafN_3542_D;
  input [63:0] base1_124_3685_D;
  input [63:0] leafvec124_3684_D;
  input [63:0] base0_118_3681_D;
  input [63:0] vec118_3676_D;
  input [63:0] base0_112_3673_D;
  input [63:0] vec112_3668_D;
  input [63:0] base0_106_3665_D;
  input [63:0] vec106_3660_D;
  input [63:0] base0_100_3657_D;
  input [63:0] vec100_3652_D;
  input [63:0] base0_94_3649_D;
  input [63:0] vec94_3644_D;
  input [63:0] base0_88_3641_D;
  input [63:0] vec88_3636_D;
  input [63:0] base0_82_3633_D;
  input [63:0] vec82_3628_D;
  input [63:0] base0_76_3625_D;
  input [63:0] vec76_3620_D;
  input [63:0] base0_70_3617_D;
  input [63:0] vec70_3612_D;
  input [63:0] base0_64_3609_D;
  input [63:0] vec64_3604_D;
  input [63:0] ip2_3602_D;
  input [63:0] base0_58_3600_D;
  input [63:0] vec58_3595_D;
  input [63:0] base0_52_3592_D;
  input [63:0] vec52_3587_D;
  input [63:0] base0_46_3584_D;
  input [63:0] vec46_3579_D;
  input [63:0] base0_40_3576_D;
  input [63:0] vec40_3571_D;
  input [63:0] base0_34_3568_D;
  input [63:0] vec34_3563_D;
  input [63:0] base0_28_3560_D;
  input [63:0] vec28_3555_D;
  input [63:0] base0_22_3552_D;
  input [63:0] vec22_3547_D;
  input [63:0] base0_16_3544_D;
  input [63:0] vec16_3538_D;
  input [63:0] dirC_3532_D;
  input [63:0] ip1_3530_D;
  //OUT
  output [7:0] R13573;
  //WIRES
  wire [7:0] R13573;
  wire [7:0] R13572;
  wire [7:0] R13571;
  wire [7:0] R13570;
  wire [7:0] R13569;
  wire [7:0] R13568;
  wire [7:0] R13567;
  wire [7:0] R13566;
  wire [63:0] R13565;
  wire [63:0] R13564;
  wire [63:0] R13563;
  wire [7:0] R13562;
  wire [7:0] R13561;
  wire [7:0] R13560;
  wire [7:0] R13559;
  wire [7:0] R13558;
  wire [7:0] R13557;
  wire [7:0] R13556;
  wire [7:0] R13555;
  wire [7:0] R13554;
  wire [7:0] R13553;
  wire [7:0] R13552;
  wire [31:0] R13551;
  wire [31:0] R13550;
  wire [63:0] R13549;
  wire [63:0] R13548;
  wire [63:0] R13547;
  wire [63:0] R13546;
  wire [63:0] R13545;
  wire [63:0] R13544;
  wire [63:0] R13543;
  wire [63:0] R13542;
  wire [7:0] R13541;
  wire [7:0] R13540;
  wire [7:0] R13539;
  wire [7:0] R13538;
  wire [7:0] R13537;
  wire [7:0] R13536;
  wire [7:0] R13535;
  wire [7:0] R13534;
  wire [7:0] R13533;
  wire [31:0] R13532;
  wire [31:0] R13531;
  wire [31:0] R13530;
  wire [31:0] R13529;
  wire [31:0] R13528;
  wire [31:0] R13527;
  wire [31:0] R13526;
  wire [31:0] R13525;
  wire [63:0] R13524;
  wire [63:0] R13523;
  wire [63:0] R13522;
  wire [63:0] R13521;
  wire [63:0] R13520;
  wire [63:0] R13519;
  wire [63:0] R13518;
  wire [63:0] R13517;
  wire [63:0] R13516;
  wire [63:0] R13515;
  wire [63:0] R13514;
  wire [31:0] R13513;
  wire [31:0] R13512;
  wire [31:0] R13511;
  wire [31:0] R13510;
  wire [31:0] R13509;
  wire [31:0] R13508;
  wire [31:0] R13507;
  wire [31:0] R13506;
  wire [31:0] R13505;
  wire [31:0] R13504;
  wire [31:0] R13503;
  wire [63:0] R13502;
  wire [63:0] R13501;
  wire [63:0] R13500;
  wire [63:0] R13499;
  wire [63:0] R13498;
  wire [63:0] R13497;
  wire [63:0] R13496;
  wire [63:0] R13495;
  wire [63:0] R13494;
  wire [63:0] R13493;
  wire [63:0] R13492;
  wire [63:0] R13491;
  wire [31:0] R13490;
  wire [31:0] R13489;
  wire [31:0] R13488;
  wire [31:0] R13487;
  wire [31:0] R13486;
  wire [31:0] R13485;
  wire [31:0] R13484;
  wire [31:0] R13483;
  wire [63:0] R13482;
  wire [63:0] R13481;
  wire [63:0] R13480;
  wire [63:0] R13479;
  wire [63:0] R13478;
  wire [63:0] R13477;
  wire [63:0] R13476;
  wire [63:0] R13475;
  wire [63:0] R13474;
  wire [63:0] R13473;
  wire [63:0] R13472;
  wire [63:0] R13471;
  wire [63:0] R13470;
  wire [63:0] R13469;
  wire [63:0] R13468;
  wire [63:0] R13467;
  wire [63:0] R13466;
  wire [63:0] R13465;
  wire [63:0] R13464;
  wire [63:0] R13463;
  wire [63:0] R13462;
  wire [63:0] R13461;
  wire [63:0] R13460;
  wire [63:0] R13459;
  wire [63:0] R13458;
  wire [63:0] R13457;
  wire [63:0] R13456;
  wire [63:0] R13455;
  wire [63:0] R13454;
  wire [31:0] R13453;
  wire [31:0] R13452;
  wire [31:0] R13451;
  wire [31:0] R13450;
  wire [31:0] R13449;
  wire [31:0] R13448;
  wire [31:0] R13447;
  wire [31:0] R13446;
  wire [31:0] R13445;
  wire [63:0] R13444;
  wire [63:0] R13443;
  wire [63:0] R13442;
  wire [63:0] R13441;
  wire [63:0] R13440;
  wire [63:0] R13439;
  wire [63:0] R13438;
  wire [63:0] R13437;
  wire [63:0] R13436;
  wire [63:0] R13435;
  wire [63:0] R13434;
  wire [63:0] R13433;
  wire [63:0] R13432;
  wire [63:0] R13431;
  wire [63:0] R13430;
  wire [63:0] R13429;
  wire [63:0] R13428;
  wire [63:0] R13427;
  wire [63:0] R13426;
  wire [63:0] R13425;
  wire [63:0] R13424;
  wire [63:0] R13423;
  wire [63:0] R13422;
  wire [63:0] R13421;
  wire [63:0] R13420;
  wire [63:0] R13419;
  wire [63:0] R13418;
  wire [63:0] R13417;
  wire [63:0] R13416;
  wire [63:0] R13415;
  wire [63:0] R13414;
  wire [63:0] R13413;
  wire [63:0] R13412;
  wire [63:0] R13411;
  wire [63:0] R13410;
  wire [63:0] R13409;
  wire [63:0] R13408;
  wire [63:0] R13407;
  wire [63:0] R13406;
  wire [63:0] R13405;
  wire [63:0] R13404;
  wire [63:0] R13403;
  wire [63:0] R13402;
  wire [63:0] R13401;
  wire [63:0] R13400;
  wire [63:0] R13399;
  wire [63:0] R13398;
  wire [63:0] R13397;
  wire [63:0] R13396;
  wire [63:0] R13395;
  wire [63:0] R13394;
  wire [63:0] R13393;
  wire [63:0] R13392;
  wire [63:0] R13391;
  wire [63:0] R13390;
  wire [63:0] R13389;
  wire [63:0] R13388;
  wire [63:0] R13387;
  wire [63:0] R13386;
  wire [63:0] R13385;
  wire [63:0] R13384;
  wire [63:0] R13383;
  wire [63:0] R13382;
  wire [63:0] R13381;
  wire [63:0] R13380;
  wire [63:0] R13379;
  wire [63:0] R13378;
  wire [63:0] R13377;
  wire [63:0] R13376;
  wire [63:0] R13375;
  wire [63:0] R13374;
  wire [63:0] R13373;
  wire [63:0] R13372;
  wire [63:0] R13371;
  wire [63:0] R13370;
  wire [63:0] R13369;
  wire [63:0] R13368;
  wire [63:0] R13367;
  wire [63:0] R13366;
  wire [63:0] R13365;
  wire [63:0] R13364;
  wire [63:0] R13363;
  wire [63:0] R13362;
  wire [63:0] R13361;
  wire [63:0] R13360;
  wire [63:0] R13359;
  wire [63:0] R13358;
  wire [63:0] R13357;
  wire [63:0] R13356;
  wire [63:0] R13355;
  wire [63:0] R13354;
  wire [63:0] R13353;
  wire [63:0] R13352;
  wire [63:0] R13351;
  wire [63:0] R13350;
  wire [63:0] R13349;
  wire [63:0] R13348;
  wire [63:0] R13347;
  wire [63:0] R13346;
  wire [63:0] R13345;
  wire [63:0] R13344;
  wire [63:0] R13343;
  wire [63:0] R13342;
  wire [63:0] R13341;
  wire [63:0] R13340;
  wire [63:0] R13339;
  wire [63:0] R13338;
  wire [63:0] R13337;
  wire [63:0] R13336;
  wire [63:0] R13335;
  wire [63:0] R13334;
  wire [63:0] R13333;
  wire [63:0] R13332;
  wire [63:0] R13331;
  wire [63:0] R13330;
  wire [63:0] R13329;
  wire [63:0] R13328;
  wire [63:0] R13327;
  wire [63:0] R13326;
  wire [63:0] R13325;
  wire [63:0] R13324;
  wire [63:0] R13323;
  wire [63:0] R13322;
  wire [63:0] R13321;
  wire [63:0] R13320;
  wire [63:0] R13319;
  wire [63:0] R13318;
  wire [63:0] R13317;
  wire [63:0] R13316;
  wire [63:0] R13315;
  wire [63:0] R13314;
  wire [63:0] R13313;
  wire [63:0] R13312;
  wire [63:0] R13311;
  wire [63:0] R13310;
  wire [63:0] R13309;
  wire [63:0] R13308;
  wire [63:0] R13307;
  wire [63:0] R13306;
  wire [63:0] R13305;
  wire [63:0] R13304;
  wire [63:0] R13303;
  wire [63:0] R13302;
  wire [63:0] R13301;
  wire [63:0] R13300;
  wire [63:0] R13299;
  wire [63:0] R13298;
  wire [63:0] R13297;
  wire [63:0] R13296;
  wire [63:0] R13295;
  wire [63:0] R13294;
  wire [63:0] R13293;
  wire [63:0] R13292;
  wire [63:0] R13291;
  wire [63:0] R13290;
  wire [63:0] R13289;
  wire [63:0] R13288;
  wire [63:0] R13287;
  wire [63:0] R13286;
  wire [63:0] R13285;
  wire [63:0] R13284;
  wire [63:0] R13283;
  wire [63:0] R13282;
  wire [63:0] R13281;
  wire [63:0] R13280;
  wire [63:0] R13279;
  wire [63:0] R13278;
  wire [63:0] R13277;
  wire [63:0] R13276;
  wire [63:0] R13275;
  wire [63:0] R13274;
  wire [63:0] R13273;
  wire [63:0] R13272;
  wire [63:0] R13271;
  wire [63:0] R13270;
  wire [63:0] R13269;
  wire [63:0] R13268;
  wire [63:0] R13267;
  wire [63:0] R13266;
  wire [63:0] R13265;
  wire [63:0] R13264;
  wire [63:0] R13263;
  wire [63:0] R13262;
  wire [63:0] R13261;
  wire [63:0] R13260;
  wire [63:0] R13259;
  wire [63:0] R13258;
  wire [63:0] R13257;
  wire [63:0] R13256;
  wire [63:0] R13255;
  wire [63:0] R13254;
  wire [63:0] R13253;
  wire [63:0] R13252;
  wire [63:0] R13251;
  wire [63:0] R13250;
  wire [63:0] R13249;
  wire [63:0] R13248;
  wire [63:0] R13247;
  wire [63:0] R13246;
  wire [63:0] R13245;
  wire [63:0] R13244;
  wire [63:0] R13243;
  wire [63:0] R13242;
  wire [63:0] R13241;
  wire [63:0] R13240;
  wire [63:0] R13239;
  wire [63:0] R13238;
  wire [63:0] R13237;
  wire [63:0] R13236;
  wire [63:0] R13235;
  wire [63:0] R13234;
  wire [63:0] R13233;
  wire [63:0] R13232;
  wire [63:0] R13231;
  wire [63:0] R13230;
  wire [63:0] R13229;
  wire [63:0] R13228;
  wire [63:0] R13227;
  wire [63:0] R13226;
  wire [63:0] R13225;
  wire [63:0] R13224;
  wire [63:0] R13223;
  wire [63:0] R13222;
  wire [63:0] R13221;
  wire [63:0] R13220;
  wire [63:0] R13219;
  wire [63:0] R13218;
  wire [63:0] R13217;
  wire [63:0] R13216;
  wire [63:0] R13215;
  wire [63:0] R13214;
  wire [63:0] R13213;
  wire [63:0] R13212;
  wire [63:0] R13211;
  wire [63:0] R13210;
  wire [63:0] R13209;
  wire [63:0] R13208;
  wire [63:0] R13207;
  wire [63:0] R13206;
  wire [63:0] R13205;
  wire [63:0] R13204;
  wire [63:0] R13203;
  wire [63:0] R13202;
  wire [63:0] R13201;
  wire [63:0] R13200;
  wire [63:0] R13199;
  wire [63:0] R13198;
  wire [63:0] R13197;
  wire [63:0] R13196;
  wire [63:0] R13195;
  wire [63:0] R13194;
  wire [63:0] R13193;
  wire [63:0] R13192;
  wire [63:0] R13191;
  wire [63:0] R13190;
  wire [63:0] R13189;
  wire [63:0] R13188;
  wire [63:0] R13187;
  wire [63:0] R13186;
  wire [63:0] R13185;
  wire [63:0] R13184;
  wire [63:0] R13183;
  wire [63:0] R13182;
  wire [63:0] R13181;
  wire [63:0] R13180;
  wire [63:0] R13179;
  wire [63:0] R13178;
  wire [63:0] R13177;
  wire [63:0] R13176;
  wire [63:0] R13175;
  wire [63:0] R13174;
  wire [63:0] R13173;
  wire [63:0] R13172;
  wire [63:0] R13171;
  wire [63:0] R13170;
  wire [63:0] R13169;
  wire [63:0] R13168;
  wire [63:0] R13167;
  wire [63:0] R13166;
  wire [63:0] R13165;
  wire [63:0] R13164;
  wire [63:0] R13163;
  wire [63:0] R13162;
  wire [63:0] R13161;
  wire [63:0] R13160;
  wire [63:0] R13159;
  wire [63:0] R13158;
  wire [63:0] R13157;
  wire [63:0] R13156;
  wire [63:0] R13155;
  wire [63:0] R13154;
  wire [63:0] R13153;
  wire [63:0] R13152;
  wire [63:0] R13151;
  wire [63:0] R13150;
  wire [63:0] R13149;
  wire [63:0] R13148;
  wire [63:0] R13147;
  wire [63:0] R13146;
  wire [63:0] R13145;
  wire [63:0] R13144;
  wire [63:0] R13143;
  wire [63:0] R13142;
  wire [63:0] R13141;
  wire [63:0] R13140;
  wire [63:0] R13139;
  wire [63:0] R13138;
  wire [63:0] R13137;
  wire [63:0] R13136;
  wire [63:0] R13135;
  wire [63:0] R13134;
  wire [63:0] R13133;
  wire [63:0] R13132;
  wire [63:0] R13131;
  wire [63:0] R13130;
  wire [63:0] R13129;
  wire [63:0] R13128;
  wire [63:0] R13127;
  wire [63:0] R13126;
  wire [63:0] R13125;
  wire [63:0] R13124;
  wire [63:0] R13123;
  wire [63:0] R13122;
  wire [63:0] R13121;
  wire [63:0] R13120;
  wire [63:0] R13119;
  wire [63:0] R13118;
  wire [63:0] R13117;
  wire [63:0] R13116;
  wire [63:0] R13115;
  wire [63:0] R13114;
  wire [63:0] R13113;
  wire [63:0] R13112;
  wire [63:0] R13111;
  wire [63:0] R13110;
  wire [63:0] R13109;
  wire [63:0] R13108;
  wire [63:0] R13107;
  wire [63:0] R13106;
  wire [63:0] R13105;
  wire [63:0] R13104;
  wire [63:0] R13103;
  wire [63:0] R13102;
  wire [63:0] R13101;
  wire [63:0] R13100;
  wire [63:0] R13099;
  wire [63:0] R13098;
  wire [63:0] R13097;
  wire [63:0] R13096;
  wire [63:0] R13095;
  wire [63:0] R13094;
  wire [63:0] R13093;
  wire [63:0] R13092;
  wire [63:0] R13091;
  wire [63:0] R13090;
  wire [63:0] R13089;
  wire [63:0] R13088;
  wire [63:0] R13087;
  wire [63:0] R13086;
  wire [63:0] R13085;
  wire [63:0] R13084;
  wire [63:0] R13083;
  wire [63:0] R13082;
  wire [63:0] R13081;
  wire [63:0] R13080;
  wire [63:0] R13079;
  wire [63:0] R13078;
  wire [63:0] R13077;
  wire [63:0] R13076;
  wire [63:0] R13075;
  wire [63:0] R13074;
  wire [63:0] R13073;
  wire [63:0] R13072;
  wire [63:0] R13071;
  wire [63:0] R13070;
  wire [63:0] R13069;
  wire [63:0] R13068;
  wire [63:0] R13067;
  wire [63:0] R13066;
  wire [63:0] R13065;
  wire [63:0] R13064;
  wire [63:0] R13063;
  wire [63:0] R13062;
  wire [63:0] R13061;
  wire [63:0] R13060;
  wire [63:0] R13059;
  wire [63:0] R13058;
  wire [63:0] R13057;
  wire [63:0] R13056;
  wire [63:0] R13055;
  wire [63:0] R13054;
  wire [63:0] R13053;
  wire [63:0] R13052;
  wire [63:0] R13051;
  wire [63:0] R13050;
  wire [63:0] R13049;
  wire [63:0] R13048;
  wire [63:0] R13047;
  wire [63:0] R13046;
  wire [63:0] R13045;
  wire [63:0] R13044;
  wire [63:0] R13043;
  wire [63:0] R13042;
  wire [63:0] R13041;
  wire [63:0] R13040;
  wire [63:0] R13039;
  wire [63:0] R13038;
  wire [63:0] R13037;
  wire [63:0] R13036;
  wire [63:0] R13035;
  wire [63:0] R13034;
  wire [63:0] R13033;
  wire [63:0] R13032;
  wire [63:0] R13031;
  wire [63:0] R13030;
  wire [63:0] R13029;
  wire [63:0] R13028;
  wire [63:0] R13027;
  wire [63:0] R13026;
  wire [63:0] R13025;
  wire [63:0] R13024;
  wire [63:0] R13023;
  wire [63:0] R13022;
  wire [63:0] R13021;
  wire [63:0] R13020;
  wire [63:0] R13019;
  wire [63:0] R13018;
  wire [63:0] R13017;
  wire [63:0] R13016;
  wire [63:0] R13015;
  wire [63:0] R13014;
  wire [63:0] R13013;
  wire [63:0] R13012;
  wire [63:0] R13011;
  wire [63:0] R13010;
  wire [63:0] R13009;
  wire [63:0] R13008;
  wire [63:0] R13007;
  wire [63:0] R13006;
  wire [63:0] R13005;
  wire [63:0] R13004;
  wire [63:0] R13003;
  wire [63:0] R13002;
  wire [63:0] R13001;
  wire [63:0] R13000;
  wire [63:0] R12999;
  wire [63:0] R12998;
  wire [63:0] R12997;
  wire [63:0] R12996;
  wire [63:0] R12995;
  wire [63:0] R12994;
  wire [63:0] R12993;
  wire [63:0] R12992;
  wire [63:0] R12991;
  wire [63:0] R12990;
  wire [63:0] R12989;
  wire [63:0] R12988;
  wire [63:0] R12987;
  wire [63:0] R12986;
  wire [63:0] R12985;
  wire [63:0] R12984;
  wire [63:0] R12983;
  wire [63:0] R12982;
  wire [63:0] R12981;
  wire [63:0] R12980;
  wire [63:0] R12979;
  wire [63:0] R12978;
  wire [63:0] R12977;
  wire [63:0] R12976;
  wire [63:0] R12975;
  wire [63:0] R12974;
  wire [63:0] R12973;
  wire [63:0] R12972;
  wire [63:0] R12971;
  wire [63:0] R12970;
  wire [63:0] R12969;
  wire [63:0] R12968;
  wire [63:0] R12967;
  wire [63:0] R12966;
  wire [63:0] R12965;
  wire [63:0] R12964;
  wire [63:0] R12963;
  wire [63:0] R12962;
  wire [63:0] R12961;
  wire [63:0] R12960;
  wire [63:0] R12959;
  wire [63:0] R12958;
  wire [63:0] R12957;
  wire [63:0] R12956;
  wire [63:0] R12955;
  wire [63:0] R12954;
  wire [63:0] R12953;
  wire [63:0] R12952;
  wire [63:0] R12951;
  wire [63:0] R12950;
  wire [63:0] R12949;
  wire [63:0] R12948;
  wire [63:0] R12947;
  wire [63:0] R12946;
  wire [63:0] R12945;
  wire [63:0] R12944;
  wire [63:0] R12943;
  wire [63:0] R12942;
  wire [63:0] R12941;
  wire [63:0] R12940;
  wire [63:0] R12939;
  wire [63:0] R12938;
  wire [63:0] R12937;
  wire [63:0] R12936;
  wire [63:0] R12935;
  wire [63:0] R12934;
  wire [63:0] R12933;
  wire [63:0] R12932;
  wire [63:0] R12931;
  wire [63:0] R12930;
  wire [63:0] R12929;
  wire [63:0] R12928;
  wire [63:0] R12927;
  wire [63:0] R12926;
  wire [63:0] R12925;
  wire [63:0] R12924;
  wire [63:0] R12923;
  wire [63:0] R12922;
  wire [63:0] R12921;
  wire [63:0] R12920;
  wire [63:0] R12919;
  wire [63:0] R12918;
  wire [63:0] R12917;
  wire [63:0] R12916;
  wire [63:0] R12915;
  wire [63:0] R12914;
  wire [63:0] R12913;
  wire [63:0] R12912;
  wire [63:0] R12911;
  wire [63:0] R12910;
  wire [63:0] R12909;
  wire [63:0] R12908;
  wire [63:0] R12907;
  wire [63:0] R12906;
  wire [63:0] R12905;
  wire [63:0] R12904;
  wire [63:0] R12903;
  wire [63:0] R12902;
  wire [63:0] R12901;
  wire [63:0] R12900;
  wire [63:0] R12899;
  wire [63:0] R12898;
  wire [63:0] R12897;
  wire [63:0] R12896;
  wire [63:0] R12895;
  wire [63:0] R12894;
  wire [63:0] R12893;
  wire [63:0] R12892;
  wire [63:0] R12891;
  wire [63:0] R12890;
  wire [63:0] R12889;
  wire [63:0] R12888;
  wire [63:0] R12887;
  wire [63:0] R12886;
  wire [63:0] R12885;
  wire [63:0] R12884;
  wire [63:0] R12883;
  wire [63:0] R12882;
  wire [63:0] R12881;
  wire [63:0] R12880;
  wire [63:0] R12879;
  wire [63:0] R12878;
  wire [63:0] R12877;
  wire [63:0] R12876;
  wire [63:0] R12875;
  wire [63:0] R12874;
  wire [63:0] R12873;
  wire [63:0] R12872;
  wire [63:0] R12871;
  wire [63:0] R12870;
  wire [63:0] R12869;
  wire [63:0] R12868;
  wire [63:0] R12867;
  wire [63:0] R12866;
  wire [63:0] R12865;
  wire [63:0] R12864;
  wire [63:0] R12863;
  wire [63:0] R12862;
  wire [63:0] R12861;
  wire [63:0] R12860;
  wire [63:0] R12859;
  wire [63:0] R12858;
  wire [63:0] R12857;
  wire [63:0] R12856;
  wire [63:0] R12855;
  wire [63:0] R12854;
  wire [63:0] R12853;
  wire [63:0] R12852;
  wire [63:0] R12851;
  wire [63:0] R12850;
  wire [63:0] R12849;
  wire [63:0] R12848;
  wire [63:0] R12847;
  wire [63:0] R12846;
  wire [63:0] R12845;
  wire [63:0] R12844;
  wire [63:0] R12843;
  wire [63:0] R12842;
  wire [63:0] R12841;
  wire [63:0] R12840;
  wire [63:0] R12839;
  wire [63:0] R12838;
  wire [63:0] R12837;
  wire [63:0] R12836;
  wire [63:0] R12835;
  wire [63:0] R12834;
  wire [63:0] R12833;
  wire [63:0] R12832;
  wire [63:0] R12831;
  wire [63:0] R12830;
  wire [63:0] R12829;
  wire [63:0] R12828;
  wire [63:0] R12827;
  wire [63:0] R12826;
  wire [63:0] R12825;
  wire [63:0] R12824;
  wire [63:0] R12823;
  wire [63:0] R12822;
  wire [63:0] R12821;
  wire [63:0] R12820;
  wire [63:0] R12819;
  wire [63:0] R12818;
  wire [63:0] R12817;
  wire [63:0] R12816;
  wire [63:0] R12815;
  wire [63:0] R12814;
  wire [63:0] R12813;
  wire [63:0] R12812;
  wire [63:0] R12811;
  wire [63:0] R12810;
  wire [63:0] R12809;
  wire [63:0] R12808;
  wire [63:0] R12807;
  wire [63:0] R12806;
  wire [63:0] R12805;
  wire [63:0] R12804;
  wire [63:0] R12803;
  wire [63:0] R12802;
  wire [63:0] R12801;
  wire [63:0] R12800;
  wire [63:0] R12799;
  wire [63:0] R12798;
  wire [63:0] R12797;
  wire [63:0] R12796;
  wire [63:0] R12795;
  wire [63:0] R12794;
  wire [63:0] R12793;
  wire [63:0] R12792;
  wire [63:0] R12791;
  wire [63:0] R12790;
  wire [63:0] R12789;
  wire [63:0] R12788;
  wire [63:0] R12787;
  wire [63:0] R12786;
  wire [63:0] R12785;
  wire [63:0] R12784;
  wire [63:0] R12783;
  wire [63:0] R12782;
  wire [63:0] R12781;
  wire [63:0] R12780;
  wire [0:0] R12779;
  wire [0:0] R12778;
  wire [0:0] R12777;
  wire [0:0] R12776;
  wire [0:0] R12775;
  wire [0:0] R12774;
  wire [0:0] R12773;
  wire [0:0] R12772;
  wire [0:0] R12771;
  wire [0:0] R12770;
  wire [0:0] R12769;
  wire [0:0] R12768;
  wire [0:0] R12767;
  wire [0:0] R12766;
  wire [0:0] R12765;
  wire [0:0] R12764;
  wire [0:0] R12763;
  wire [0:0] R12762;
  wire [0:0] R12761;
  wire [0:0] R12760;
  wire [0:0] R12759;
  wire [0:0] R12758;
  wire [63:0] R12757;
  wire [63:0] R12756;
  wire [63:0] R12755;
  wire [63:0] R12754;
  wire [63:0] R12753;
  wire [63:0] R12752;
  wire [63:0] R12751;
  wire [63:0] R12750;
  wire [63:0] R12749;
  wire [63:0] R12748;
  wire [63:0] R12747;
  wire [63:0] R12746;
  wire [63:0] R12745;
  wire [63:0] R12744;
  wire [63:0] R12743;
  wire [63:0] R12742;
  wire [63:0] R12741;
  wire [63:0] R12740;
  wire [63:0] R12739;
  wire [63:0] R12738;
  wire [63:0] R12737;
  wire [63:0] R12736;
  wire [63:0] R12735;
  wire [63:0] R12734;
  wire [63:0] R12733;
  wire [63:0] R12732;
  wire [63:0] R12731;
  wire [63:0] R12730;
  wire [63:0] R12729;
  wire [63:0] R12728;
  wire [63:0] R12727;
  wire [63:0] R12726;
  wire [63:0] R12725;
  wire [63:0] R12724;
  wire [63:0] R12723;
  wire [63:0] R12722;
  wire [63:0] R12721;
  wire [63:0] R12720;
  wire [63:0] R12719;
  wire [63:0] R12718;
  wire [63:0] R12717;
  wire [63:0] R12716;
  wire [63:0] R12715;
  wire [63:0] R12714;
  wire [63:0] R12713;
  wire [63:0] R12712;
  wire [63:0] R12711;
  wire [63:0] R12710;
  wire [63:0] R12709;
  wire [63:0] R12708;
  wire [63:0] R12707;
  wire [63:0] R12706;
  wire [63:0] R12705;
  wire [63:0] R12704;
  wire [63:0] R12703;
  wire [63:0] R12702;
  wire [63:0] R12701;
  wire [63:0] R12700;
  wire [63:0] R12699;
  wire [63:0] R12698;
  wire [63:0] R12697;
  wire [63:0] R12696;
  wire [63:0] R12695;
  wire [63:0] R12694;
  wire [63:0] R12693;
  wire [63:0] R12692;
  wire [63:0] R12691;
  wire [63:0] R12690;
  wire [63:0] R12689;
  wire [63:0] R12688;
  wire [63:0] R12687;
  wire [63:0] R12686;
  wire [63:0] R12685;
  wire [63:0] R12684;
  wire [63:0] R12683;
  wire [63:0] R12682;
  wire [63:0] R12681;
  wire [63:0] R12680;
  wire [63:0] R12679;
  wire [63:0] R12678;
  wire [63:0] R12677;
  wire [63:0] R12676;
  wire [63:0] R12675;
  wire [63:0] R12674;
  wire [63:0] R12673;
  wire [63:0] R12672;
  wire [63:0] R12671;
  wire [63:0] R12670;
  wire [63:0] R12669;
  wire [63:0] R12668;
  wire [63:0] R12667;
  wire [63:0] R12666;
  wire [63:0] R12665;
  wire [63:0] R12664;
  wire [63:0] R12663;
  wire [63:0] R12662;
  wire [63:0] R12661;
  wire [63:0] R12660;
  wire [63:0] R12659;
  wire [63:0] R12658;
  wire [63:0] R12657;
  wire [63:0] R12656;
  wire [63:0] R12655;
  wire [63:0] R12654;
  wire [63:0] R12653;
  wire [63:0] R12652;
  wire [63:0] R12651;
  wire [63:0] R12650;
  wire [63:0] R12649;
  wire [63:0] R12648;
  wire [63:0] R12647;
  wire [63:0] R12646;
  wire [63:0] R12645;
  wire [63:0] R12644;
  wire [63:0] R12643;
  wire [63:0] R12642;
  wire [63:0] R12641;
  wire [63:0] R12640;
  wire [63:0] R12639;
  wire [63:0] R12638;
  wire [63:0] R12637;
  wire [63:0] R12636;
  wire [63:0] R12635;
  wire [63:0] R12634;
  wire [63:0] R12633;
  wire [63:0] R12632;
  wire [63:0] R12631;
  wire [63:0] R12630;
  wire [63:0] R12629;
  wire [63:0] R12628;
  wire [63:0] R12627;
  wire [63:0] R12626;
  wire [63:0] R12625;
  wire [63:0] R12624;
  wire [63:0] R12623;
  wire [63:0] R12622;
  wire [63:0] R12621;
  wire [63:0] R12620;
  wire [63:0] R12619;
  wire [63:0] R12618;
  wire [63:0] R12617;
  wire [63:0] R12616;
  wire [63:0] R12615;
  wire [63:0] R12614;
  wire [63:0] R12613;
  wire [63:0] R12612;
  wire [63:0] R12611;
  wire [63:0] R12610;
  wire [63:0] R12609;
  wire [63:0] R12608;
  wire [63:0] R12607;
  wire [0:0] R12606;
  wire [0:0] R12605;
  wire [0:0] R12604;
  wire [0:0] R12603;
  wire [0:0] R12602;
  wire [0:0] R12601;
  wire [0:0] R12600;
  wire [0:0] R12599;
  wire [0:0] R12598;
  wire [0:0] R12597;
  wire [0:0] R12596;
  wire [0:0] R12595;
  wire [0:0] R12594;
  wire [0:0] R12593;
  wire [0:0] R12592;
  wire [0:0] R12591;
  wire [0:0] R12590;
  wire [0:0] R12589;
  wire [0:0] R12588;
  wire [0:0] R12587;
  wire [0:0] R12586;
  wire [0:0] R12585;
  wire [0:0] R12584;
  wire [0:0] R12583;
  wire [0:0] R12582;
  wire [0:0] R12581;
  wire [0:0] R12580;
  wire [0:0] R12579;
  wire [0:0] R12578;
  wire [0:0] R12577;
  wire [0:0] R12576;
  wire [0:0] R12575;
  wire [0:0] R12574;
  wire [0:0] R12573;
  wire [0:0] R12572;
  wire [0:0] R12571;
  wire [0:0] R12570;
  wire [0:0] R12569;
  wire [0:0] R12568;
  wire [0:0] R12567;
  wire [0:0] R12566;
  wire [0:0] R12565;
  wire [0:0] R12564;
  wire [0:0] R12563;
  wire [0:0] R12562;
  wire [0:0] R12561;
  wire [0:0] R12560;
  wire [0:0] R12559;
  wire [0:0] R12558;
  wire [0:0] R12557;
  wire [0:0] R12556;
  wire [0:0] R12555;
  wire [0:0] R12554;
  wire [0:0] R12553;
  wire [0:0] R12552;
  wire [0:0] R12551;
  wire [0:0] R12550;
  wire [0:0] R12549;
  wire [0:0] R12548;
  wire [0:0] R12547;
  wire [0:0] R12546;
  wire [0:0] R12545;
  wire [0:0] R12544;
  wire [0:0] R12543;
  wire [0:0] R12542;
  wire [0:0] R12541;
  wire [0:0] R12540;
  wire [0:0] R12539;
  wire [0:0] R12538;
  wire [0:0] R12537;
  wire [0:0] R12536;
  wire [0:0] R12535;
  wire [0:0] R12534;
  wire [0:0] R12533;
  wire [0:0] R12532;
  wire [0:0] R12531;
  wire [0:0] R12530;
  wire [0:0] R12529;
  wire [0:0] R12528;
  wire [0:0] R12527;
  wire [0:0] R12526;
  wire [0:0] R12525;
  wire [0:0] R12524;
  wire [0:0] R12523;
  wire [0:0] R12522;
  wire [0:0] R12521;
  wire [0:0] R12520;
  wire [0:0] R12519;
  wire [63:0] R12518;
  wire [63:0] R12517;
  wire [63:0] R12516;
  wire [63:0] R12515;
  wire [63:0] R12514;
  wire [63:0] R12513;
  wire [63:0] R12512;
  wire [63:0] R12511;
  wire [63:0] R12510;
  wire [63:0] R12509;
  wire [63:0] R12508;
  wire [63:0] R12507;
  wire [63:0] R12506;
  wire [63:0] R12505;
  wire [63:0] R12504;
  wire [63:0] R12503;
  wire [63:0] R12502;
  wire [63:0] R12501;
  wire [63:0] R12500;
  wire [63:0] R12499;
  wire [63:0] R12498;
  wire [63:0] R12497;
  wire [63:0] R12496;
  wire [63:0] R12495;
  wire [63:0] R12494;
  wire [63:0] R12493;
  wire [63:0] R12492;
  wire [63:0] R12491;
  wire [63:0] R12490;
  wire [63:0] R12489;
  wire [63:0] R12488;
  wire [63:0] R12487;
  wire [63:0] R12486;
  wire [63:0] R12485;
  wire [63:0] R12484;
  wire [63:0] R12483;
  wire [63:0] R12482;
  wire [63:0] R12481;
  wire [63:0] R12480;
  wire [63:0] R12479;
  wire [63:0] R12478;
  wire [63:0] R12477;
  wire [63:0] R12476;
  wire [63:0] R12475;
  wire [0:0] R12474;
  wire [0:0] R12473;
  wire [0:0] R12472;
  wire [0:0] R12471;
  wire [0:0] R12470;
  wire [0:0] R12469;
  wire [0:0] R12468;
  wire [0:0] R12467;
  wire [0:0] R12466;
  wire [0:0] R12465;
  wire [0:0] R12464;
  wire [0:0] R12463;
  wire [0:0] R12462;
  wire [0:0] R12461;
  wire [0:0] R12460;
  wire [0:0] R12459;
  wire [0:0] R12458;
  wire [0:0] R12457;
  wire [0:0] R12456;
  wire [0:0] R12455;
  wire [0:0] R12454;
  wire [0:0] R12453;
  wire [0:0] R12452;
  wire [0:0] R12451;
  wire [0:0] R12450;
  wire [0:0] R12449;
  wire [0:0] R12448;
  wire [0:0] R12447;
  wire [0:0] R12446;
  wire [0:0] R12445;
  wire [0:0] R12444;
  wire [0:0] R12443;
  wire [0:0] R12442;
  wire [0:0] R12441;
  wire [0:0] R12440;
  wire [0:0] R12439;
  wire [0:0] R12438;
  wire [0:0] R12437;
  wire [0:0] R12436;
  wire [0:0] R12435;
  wire [0:0] R12434;
  wire [0:0] R12433;
  wire [0:0] R12432;
  wire [0:0] R12431;
  wire [0:0] R12430;
  wire [0:0] R12429;
  wire [0:0] R12428;
  wire [0:0] R12427;
  wire [0:0] R12426;
  wire [0:0] R12425;
  wire [0:0] R12424;
  wire [0:0] R12423;
  wire [0:0] R12422;
  wire [0:0] R12421;
  wire [0:0] R12420;
  wire [0:0] R12419;
  wire [0:0] R12418;
  wire [0:0] R12417;
  wire [0:0] R12416;
  wire [0:0] R12415;
  wire [0:0] R12414;
  wire [0:0] R12413;
  wire [0:0] R12412;
  wire [0:0] R12411;
  wire [0:0] R12410;
  wire [0:0] R12409;
  wire [0:0] R12408;
  wire [0:0] R12407;
  wire [0:0] R12406;
  wire [0:0] R12405;
  wire [0:0] R12404;
  wire [0:0] R12403;
  wire [0:0] R12402;
  wire [0:0] R12401;
  wire [0:0] R12400;
  wire [0:0] R12399;
  wire [0:0] R12398;
  wire [0:0] R12397;
  wire [0:0] R12396;
  wire [0:0] R12395;
  wire [0:0] R12394;
  wire [0:0] R12393;
  wire [0:0] R12392;
  wire [0:0] R12391;
  wire [0:0] R12390;
  wire [0:0] R12389;
  wire [0:0] R12388;
  wire [0:0] R12387;
  wire [0:0] R12386;
  wire [0:0] R12385;
  wire [0:0] R12384;
  wire [0:0] R12383;
  wire [0:0] R12382;
  wire [0:0] R12381;
  wire [0:0] R12380;
  wire [0:0] R12379;
  wire [0:0] R12378;
  wire [0:0] R12377;
  wire [0:0] R12376;
  wire [63:0] R12375;
  wire [63:0] R12374;
  wire [63:0] R12373;
  wire [63:0] R12372;
  wire [63:0] R12371;
  wire [63:0] R12370;
  wire [63:0] R12369;
  wire [63:0] R12368;
  wire [63:0] R12367;
  wire [63:0] R12366;
  wire [63:0] R12365;
  wire [31:0] R12364;
  wire [31:0] R12363;
  wire [31:0] R12362;
  wire [31:0] R12361;
  wire [63:0] R12360;
  wire [63:0] R12359;
  wire [63:0] R12358;
  wire [63:0] R12357;
  wire [63:0] R12356;
  wire [63:0] R12355;
  wire [63:0] R12354;
  wire [63:0] R12353;
  wire [63:0] R12352;
  wire [63:0] R12351;
  wire [63:0] R12350;
  wire [63:0] R12349;
  wire [63:0] R12348;
  wire [63:0] R12347;
  wire [63:0] R12346;
  wire [63:0] R12345;
  wire [63:0] R12344;
  wire [63:0] R12343;
  wire [63:0] R12342;
  wire [63:0] R12341;
  wire [63:0] R12340;
  wire [63:0] R12339;
  wire [63:0] R12338;
  wire [63:0] R12337;
  wire [63:0] R12336;
  wire [63:0] R12335;
  wire [63:0] R12334;
  wire [63:0] R12333;
  wire [63:0] R12332;
  wire [63:0] R12331;
  wire [63:0] R12330;
  wire [63:0] R12329;
  wire [63:0] R12328;
  wire [63:0] R12327;
  wire [63:0] R12326;
  wire [63:0] R12325;
  wire [63:0] R12324;
  wire [63:0] R12323;
  wire [63:0] R12322;
  wire [63:0] R12321;
  wire [63:0] R12320;
  wire [63:0] R12319;
  wire [63:0] R12318;
  wire [63:0] R12317;
  wire [63:0] R12316;
  wire [63:0] R12315;
  wire [63:0] R12314;
  wire [63:0] R12313;
  wire [63:0] R12312;
  wire [63:0] R12311;
  wire [63:0] R12310;
  wire [63:0] R12309;
  wire [63:0] R12308;
  wire [63:0] R12307;
  wire [63:0] R12306;
  wire [63:0] R12305;
  wire [31:0] R12304;
  wire [31:0] R12303;
  wire [31:0] R12302;
  wire [31:0] R12301;
  wire [31:0] R12300;
  wire [31:0] R12299;
  wire [31:0] R12298;
  wire [31:0] R12297;
  wire [31:0] R12296;
  wire [31:0] R12295;
  wire [63:0] R12294;
  wire [31:0] R12293;
  wire [63:0] R12292;
  wire [63:0] R12291;
  wire [63:0] R12290;
  wire [63:0] R12289;
  wire [63:0] R12288;
  wire [63:0] R12287;
  wire [63:0] R12286;
  wire [63:0] R12285;
  wire [63:0] R12284;
  wire [63:0] R12283;
  wire [63:0] R12282;
  wire [63:0] R12281;
  wire [63:0] R12280;
  wire [63:0] R12279;
  wire [63:0] R12278;
  wire [63:0] R12277;
  wire [63:0] R12276;
  wire [63:0] R12275;
  wire [63:0] R12274;
  wire [63:0] R12273;
  wire [63:0] R12272;
  wire [63:0] R12271;
  wire [63:0] R12270;
  wire [63:0] R12269;
  wire [63:0] R12268;
  wire [63:0] R12267;
  wire [63:0] R12266;
  wire [63:0] R12265;
  wire [63:0] R12264;
  wire [63:0] R12263;
  wire [63:0] R12262;
  wire [63:0] R12261;
  wire [63:0] R12260;
  wire [63:0] R12259;
  wire [63:0] R12258;
  wire [63:0] R12257;
  wire [63:0] R12256;
  wire [63:0] R12255;
  wire [63:0] R12254;
  wire [63:0] R12253;
  wire [63:0] R12252;
  wire [63:0] R12251;
  wire [63:0] R12250;
  wire [63:0] R12249;
  wire [63:0] R12248;
  wire [63:0] R12247;
  wire [0:0] R12246;
  wire [0:0] R12245;
  wire [0:0] R12244;
  wire [0:0] R12243;
  wire [0:0] R12242;
  wire [0:0] R12241;
  wire [0:0] R12240;
  wire [0:0] R12239;
  wire [0:0] R12238;
  wire [0:0] R12237;
  wire [0:0] R12236;
  wire [0:0] R12235;
  wire [0:0] R12234;
  wire [0:0] R12233;
  wire [0:0] R12232;
  wire [0:0] R12231;
  wire [0:0] R12230;
  wire [0:0] R12229;
  wire [0:0] R12228;
  wire [0:0] R12227;
  wire [0:0] R12226;
  wire [0:0] R12225;
  wire [0:0] R12224;
  wire [0:0] R12223;
  wire [63:0] R12222;
  wire [31:0] R12221;
  wire [31:0] R12220;
  wire [31:0] R12219;
  wire [31:0] R12218;
  wire [31:0] R12217;
  wire [31:0] R12216;
  wire [31:0] R12215;
  wire [31:0] R12214;
  wire [31:0] R12213;
  wire [31:0] R12212;
  wire [31:0] R12211;
  wire [31:0] R12210;
  wire [31:0] R12209;
  wire [31:0] R12208;
  wire [31:0] R12207;
  wire [31:0] R12206;
  wire [31:0] R12205;
  wire [63:0] R12204;
  wire [63:0] R12203;
  wire [63:0] R12202;
  wire [31:0] R12201;
  wire [31:0] R12200;
  wire [31:0] R12199;
  wire [31:0] R12198;
  wire [31:0] R12197;
  wire [31:0] R12196;
  wire [31:0] R12195;
  wire [31:0] R12194;
  wire [31:0] R12193;
  wire [31:0] R12192;
  wire [31:0] R12191;
  wire [31:0] R12190;
  wire [31:0] R12189;
  wire [31:0] R12188;
  wire [31:0] R12187;
  wire [31:0] R12186;
  wire [31:0] R12185;
  wire [31:0] R12184;
  wire [31:0] R12183;
  wire [31:0] R12182;
  wire [31:0] R12181;
  wire [31:0] R12180;
  wire [31:0] R12179;
  wire [63:0] R12178;
  wire [31:0] R12177;
  wire [63:0] R12176;
  wire [63:0] R12175;
  wire [63:0] R12174;
  wire [63:0] R12173;
  wire [63:0] R12172;
  wire [63:0] R12171;
  wire [63:0] R12170;
  wire [63:0] R12169;
  wire [63:0] R12168;
  wire [63:0] R12167;
  wire [63:0] R12166;
  wire [63:0] R12165;
  wire [63:0] R12164;
  wire [63:0] R12163;
  wire [63:0] R12162;
  wire [63:0] R12161;
  wire [63:0] R12160;
  wire [63:0] R12159;
  wire [63:0] R12158;
  wire [63:0] R12157;
  wire [63:0] R12156;
  wire [63:0] R12155;
  wire [63:0] R12154;
  wire [63:0] R12153;
  wire [63:0] R12152;
  wire [63:0] R12151;
  wire [63:0] R12150;
  wire [63:0] R12149;
  wire [63:0] R12148;
  wire [63:0] R12147;
  wire [63:0] R12146;
  wire [63:0] R12145;
  wire [63:0] R12144;
  wire [63:0] R12143;
  wire [63:0] R12142;
  wire [63:0] R12141;
  wire [63:0] R12140;
  wire [63:0] R12139;
  wire [63:0] R12138;
  wire [63:0] R12137;
  wire [63:0] R12136;
  wire [63:0] R12135;
  wire [63:0] R12134;
  wire [63:0] R12133;
  wire [63:0] R12132;
  wire [63:0] R12131;
  wire [0:0] R12130;
  wire [0:0] R12129;
  wire [0:0] R12128;
  wire [0:0] R12127;
  wire [0:0] R12126;
  wire [0:0] R12125;
  wire [0:0] R12124;
  wire [0:0] R12123;
  wire [0:0] R12122;
  wire [0:0] R12121;
  wire [0:0] R12120;
  wire [0:0] R12119;
  wire [0:0] R12118;
  wire [0:0] R12117;
  wire [0:0] R12116;
  wire [0:0] R12115;
  wire [0:0] R12114;
  wire [0:0] R12113;
  wire [0:0] R12112;
  wire [0:0] R12111;
  wire [0:0] R12110;
  wire [0:0] R12109;
  wire [0:0] R12108;
  wire [0:0] R12107;
  wire [0:0] R12106;
  wire [0:0] R12105;
  wire [0:0] R12104;
  wire [0:0] R12103;
  wire [0:0] R12102;
  wire [0:0] R12101;
  wire [0:0] R12100;
  wire [0:0] R12099;
  wire [0:0] R12098;
  wire [0:0] R12097;
  wire [0:0] R12096;
  wire [0:0] R12095;
  wire [0:0] R12094;
  wire [63:0] R12093;
  wire [31:0] R12092;
  wire [31:0] R12091;
  wire [31:0] R12090;
  wire [31:0] R12089;
  wire [31:0] R12088;
  wire [31:0] R12087;
  wire [31:0] R12086;
  wire [31:0] R12085;
  wire [31:0] R12084;
  wire [31:0] R12083;
  wire [31:0] R12082;
  wire [31:0] R12081;
  wire [31:0] R12080;
  wire [31:0] R12079;
  wire [31:0] R12078;
  wire [31:0] R12077;
  wire [31:0] R12076;
  wire [31:0] R12075;
  wire [31:0] R12074;
  wire [31:0] R12073;
  wire [31:0] R12072;
  wire [31:0] R12071;
  wire [31:0] R12070;
  wire [31:0] R12069;
  wire [31:0] R12068;
  wire [31:0] R12067;
  wire [31:0] R12066;
  wire [31:0] R12065;
  wire [31:0] R12064;
  wire [31:0] R12063;
  wire [63:0] R12062;
  wire [63:0] R12061;
  wire [63:0] R12060;
  wire [31:0] R12059;
  wire [31:0] R12058;
  wire [31:0] R12057;
  wire [31:0] R12056;
  wire [31:0] R12055;
  wire [31:0] R12054;
  wire [31:0] R12053;
  wire [31:0] R12052;
  wire [31:0] R12051;
  wire [31:0] R12050;
  wire [31:0] R12049;
  wire [31:0] R12048;
  wire [31:0] R12047;
  wire [31:0] R12046;
  wire [31:0] R12045;
  wire [31:0] R12044;
  wire [31:0] R12043;
  wire [31:0] R12042;
  wire [31:0] R12041;
  wire [31:0] R12040;
  wire [31:0] R12039;
  wire [31:0] R12038;
  wire [31:0] R12037;
  wire [31:0] R12036;
  wire [31:0] R12035;
  wire [31:0] R12034;
  wire [31:0] R12033;
  wire [31:0] R12032;
  wire [31:0] R12031;
  wire [31:0] R12030;
  wire [31:0] R12029;
  wire [31:0] R12028;
  wire [31:0] R12027;
  wire [31:0] R12026;
  wire [31:0] R12025;
  wire [31:0] R12024;
  wire [63:0] R12023;
  wire [31:0] R12022;
  wire [63:0] R12021;
  wire [63:0] R12020;
  wire [63:0] R12019;
  wire [63:0] R12018;
  wire [63:0] R12017;
  wire [63:0] R12016;
  wire [63:0] R12015;
  wire [63:0] R12014;
  wire [63:0] R12013;
  wire [63:0] R12012;
  wire [63:0] R12011;
  wire [63:0] R12010;
  wire [63:0] R12009;
  wire [63:0] R12008;
  wire [63:0] R12007;
  wire [63:0] R12006;
  wire [63:0] R12005;
  wire [63:0] R12004;
  wire [63:0] R12003;
  wire [63:0] R12002;
  wire [63:0] R12001;
  wire [63:0] R12000;
  wire [63:0] R11999;
  wire [63:0] R11998;
  wire [63:0] R11997;
  wire [63:0] R11996;
  wire [63:0] R11995;
  wire [63:0] R11994;
  wire [63:0] R11993;
  wire [63:0] R11992;
  wire [63:0] R11991;
  wire [63:0] R11990;
  wire [63:0] R11989;
  wire [63:0] R11988;
  wire [63:0] R11987;
  wire [63:0] R11986;
  wire [63:0] R11985;
  wire [63:0] R11984;
  wire [63:0] R11983;
  wire [63:0] R11982;
  wire [63:0] R11981;
  wire [63:0] R11980;
  wire [63:0] R11979;
  wire [63:0] R11978;
  wire [63:0] R11977;
  wire [63:0] R11976;
  wire [0:0] R11975;
  wire [0:0] R11974;
  wire [0:0] R11973;
  wire [0:0] R11972;
  wire [0:0] R11971;
  wire [0:0] R11970;
  wire [0:0] R11969;
  wire [0:0] R11968;
  wire [0:0] R11967;
  wire [0:0] R11966;
  wire [0:0] R11965;
  wire [0:0] R11964;
  wire [0:0] R11963;
  wire [0:0] R11962;
  wire [0:0] R11961;
  wire [0:0] R11960;
  wire [0:0] R11959;
  wire [0:0] R11958;
  wire [0:0] R11957;
  wire [0:0] R11956;
  wire [0:0] R11955;
  wire [0:0] R11954;
  wire [0:0] R11953;
  wire [0:0] R11952;
  wire [0:0] R11951;
  wire [0:0] R11950;
  wire [0:0] R11949;
  wire [0:0] R11948;
  wire [0:0] R11947;
  wire [0:0] R11946;
  wire [0:0] R11945;
  wire [0:0] R11944;
  wire [0:0] R11943;
  wire [0:0] R11942;
  wire [0:0] R11941;
  wire [0:0] R11940;
  wire [0:0] R11939;
  wire [0:0] R11938;
  wire [0:0] R11937;
  wire [0:0] R11936;
  wire [0:0] R11935;
  wire [0:0] R11934;
  wire [0:0] R11933;
  wire [0:0] R11932;
  wire [0:0] R11931;
  wire [0:0] R11930;
  wire [0:0] R11929;
  wire [0:0] R11928;
  wire [0:0] R11927;
  wire [0:0] R11926;
  wire [63:0] R11925;
  wire [31:0] R11924;
  wire [31:0] R11923;
  wire [31:0] R11922;
  wire [31:0] R11921;
  wire [31:0] R11920;
  wire [31:0] R11919;
  wire [31:0] R11918;
  wire [31:0] R11917;
  wire [31:0] R11916;
  wire [31:0] R11915;
  wire [31:0] R11914;
  wire [31:0] R11913;
  wire [31:0] R11912;
  wire [31:0] R11911;
  wire [31:0] R11910;
  wire [31:0] R11909;
  wire [31:0] R11908;
  wire [31:0] R11907;
  wire [31:0] R11906;
  wire [31:0] R11905;
  wire [31:0] R11904;
  wire [31:0] R11903;
  wire [31:0] R11902;
  wire [31:0] R11901;
  wire [31:0] R11900;
  wire [31:0] R11899;
  wire [31:0] R11898;
  wire [31:0] R11897;
  wire [31:0] R11896;
  wire [31:0] R11895;
  wire [31:0] R11894;
  wire [31:0] R11893;
  wire [31:0] R11892;
  wire [31:0] R11891;
  wire [31:0] R11890;
  wire [31:0] R11889;
  wire [31:0] R11888;
  wire [31:0] R11887;
  wire [31:0] R11886;
  wire [31:0] R11885;
  wire [31:0] R11884;
  wire [31:0] R11883;
  wire [31:0] R11882;
  wire [63:0] R11881;
  wire [63:0] R11880;
  wire [63:0] R11879;
  wire [31:0] R11878;
  wire [31:0] R11877;
  wire [31:0] R11876;
  wire [31:0] R11875;
  wire [31:0] R11874;
  wire [31:0] R11873;
  wire [31:0] R11872;
  wire [31:0] R11871;
  wire [31:0] R11870;
  wire [31:0] R11869;
  wire [31:0] R11868;
  wire [31:0] R11867;
  wire [31:0] R11866;
  wire [31:0] R11865;
  wire [31:0] R11864;
  wire [31:0] R11863;
  wire [31:0] R11862;
  wire [31:0] R11861;
  wire [31:0] R11860;
  wire [31:0] R11859;
  wire [31:0] R11858;
  wire [31:0] R11857;
  wire [31:0] R11856;
  wire [31:0] R11855;
  wire [31:0] R11854;
  wire [31:0] R11853;
  wire [31:0] R11852;
  wire [31:0] R11851;
  wire [31:0] R11850;
  wire [31:0] R11849;
  wire [31:0] R11848;
  wire [31:0] R11847;
  wire [31:0] R11846;
  wire [31:0] R11845;
  wire [31:0] R11844;
  wire [31:0] R11843;
  wire [31:0] R11842;
  wire [31:0] R11841;
  wire [31:0] R11840;
  wire [31:0] R11839;
  wire [31:0] R11838;
  wire [31:0] R11837;
  wire [31:0] R11836;
  wire [31:0] R11835;
  wire [31:0] R11834;
  wire [31:0] R11833;
  wire [31:0] R11832;
  wire [31:0] R11831;
  wire [31:0] R11830;
  wire [63:0] R11829;
  wire [31:0] R11828;
  wire [63:0] R11827;
  wire [63:0] R11826;
  wire [63:0] R11825;
  wire [63:0] R11824;
  wire [63:0] R11823;
  wire [63:0] R11822;
  wire [63:0] R11821;
  wire [63:0] R11820;
  wire [63:0] R11819;
  wire [63:0] R11818;
  wire [63:0] R11817;
  wire [63:0] R11816;
  wire [63:0] R11815;
  wire [63:0] R11814;
  wire [63:0] R11813;
  wire [63:0] R11812;
  wire [63:0] R11811;
  wire [63:0] R11810;
  wire [63:0] R11809;
  wire [63:0] R11808;
  wire [63:0] R11807;
  wire [63:0] R11806;
  wire [63:0] R11805;
  wire [63:0] R11804;
  wire [63:0] R11803;
  wire [63:0] R11802;
  wire [63:0] R11801;
  wire [63:0] R11800;
  wire [63:0] R11799;
  wire [63:0] R11798;
  wire [63:0] R11797;
  wire [63:0] R11796;
  wire [63:0] R11795;
  wire [63:0] R11794;
  wire [63:0] R11793;
  wire [63:0] R11792;
  wire [63:0] R11791;
  wire [63:0] R11790;
  wire [63:0] R11789;
  wire [63:0] R11788;
  wire [63:0] R11787;
  wire [63:0] R11786;
  wire [63:0] R11785;
  wire [63:0] R11784;
  wire [63:0] R11783;
  wire [63:0] R11782;
  wire [0:0] R11781;
  wire [0:0] R11780;
  wire [0:0] R11779;
  wire [0:0] R11778;
  wire [0:0] R11777;
  wire [0:0] R11776;
  wire [0:0] R11775;
  wire [0:0] R11774;
  wire [0:0] R11773;
  wire [0:0] R11772;
  wire [0:0] R11771;
  wire [0:0] R11770;
  wire [0:0] R11769;
  wire [0:0] R11768;
  wire [0:0] R11767;
  wire [0:0] R11766;
  wire [0:0] R11765;
  wire [0:0] R11764;
  wire [0:0] R11763;
  wire [0:0] R11762;
  wire [0:0] R11761;
  wire [0:0] R11760;
  wire [0:0] R11759;
  wire [0:0] R11758;
  wire [0:0] R11757;
  wire [0:0] R11756;
  wire [0:0] R11755;
  wire [0:0] R11754;
  wire [0:0] R11753;
  wire [0:0] R11752;
  wire [0:0] R11751;
  wire [0:0] R11750;
  wire [0:0] R11749;
  wire [0:0] R11748;
  wire [0:0] R11747;
  wire [0:0] R11746;
  wire [0:0] R11745;
  wire [0:0] R11744;
  wire [0:0] R11743;
  wire [0:0] R11742;
  wire [0:0] R11741;
  wire [0:0] R11740;
  wire [0:0] R11739;
  wire [0:0] R11738;
  wire [0:0] R11737;
  wire [0:0] R11736;
  wire [0:0] R11735;
  wire [0:0] R11734;
  wire [0:0] R11733;
  wire [0:0] R11732;
  wire [0:0] R11731;
  wire [0:0] R11730;
  wire [0:0] R11729;
  wire [0:0] R11728;
  wire [0:0] R11727;
  wire [0:0] R11726;
  wire [0:0] R11725;
  wire [0:0] R11724;
  wire [0:0] R11723;
  wire [0:0] R11722;
  wire [0:0] R11721;
  wire [0:0] R11720;
  wire [0:0] R11719;
  wire [63:0] R11718;
  wire [31:0] R11717;
  wire [31:0] R11716;
  wire [31:0] R11715;
  wire [31:0] R11714;
  wire [31:0] R11713;
  wire [31:0] R11712;
  wire [31:0] R11711;
  wire [31:0] R11710;
  wire [31:0] R11709;
  wire [31:0] R11708;
  wire [31:0] R11707;
  wire [31:0] R11706;
  wire [31:0] R11705;
  wire [31:0] R11704;
  wire [31:0] R11703;
  wire [31:0] R11702;
  wire [31:0] R11701;
  wire [31:0] R11700;
  wire [31:0] R11699;
  wire [31:0] R11698;
  wire [31:0] R11697;
  wire [31:0] R11696;
  wire [31:0] R11695;
  wire [31:0] R11694;
  wire [31:0] R11693;
  wire [31:0] R11692;
  wire [31:0] R11691;
  wire [31:0] R11690;
  wire [31:0] R11689;
  wire [31:0] R11688;
  wire [31:0] R11687;
  wire [31:0] R11686;
  wire [31:0] R11685;
  wire [31:0] R11684;
  wire [31:0] R11683;
  wire [31:0] R11682;
  wire [31:0] R11681;
  wire [31:0] R11680;
  wire [31:0] R11679;
  wire [31:0] R11678;
  wire [31:0] R11677;
  wire [31:0] R11676;
  wire [31:0] R11675;
  wire [31:0] R11674;
  wire [31:0] R11673;
  wire [31:0] R11672;
  wire [31:0] R11671;
  wire [31:0] R11670;
  wire [31:0] R11669;
  wire [31:0] R11668;
  wire [31:0] R11667;
  wire [31:0] R11666;
  wire [31:0] R11665;
  wire [31:0] R11664;
  wire [31:0] R11663;
  wire [31:0] R11662;
  wire [63:0] R11661;
  wire [63:0] R11660;
  wire [63:0] R11659;
  wire [31:0] R11658;
  wire [31:0] R11657;
  wire [31:0] R11656;
  wire [31:0] R11655;
  wire [31:0] R11654;
  wire [31:0] R11653;
  wire [31:0] R11652;
  wire [31:0] R11651;
  wire [31:0] R11650;
  wire [31:0] R11649;
  wire [31:0] R11648;
  wire [31:0] R11647;
  wire [31:0] R11646;
  wire [31:0] R11645;
  wire [31:0] R11644;
  wire [31:0] R11643;
  wire [31:0] R11642;
  wire [31:0] R11641;
  wire [31:0] R11640;
  wire [31:0] R11639;
  wire [31:0] R11638;
  wire [31:0] R11637;
  wire [31:0] R11636;
  wire [31:0] R11635;
  wire [31:0] R11634;
  wire [31:0] R11633;
  wire [31:0] R11632;
  wire [31:0] R11631;
  wire [31:0] R11630;
  wire [31:0] R11629;
  wire [31:0] R11628;
  wire [31:0] R11627;
  wire [31:0] R11626;
  wire [31:0] R11625;
  wire [31:0] R11624;
  wire [31:0] R11623;
  wire [31:0] R11622;
  wire [31:0] R11621;
  wire [31:0] R11620;
  wire [31:0] R11619;
  wire [31:0] R11618;
  wire [31:0] R11617;
  wire [31:0] R11616;
  wire [31:0] R11615;
  wire [31:0] R11614;
  wire [31:0] R11613;
  wire [31:0] R11612;
  wire [31:0] R11611;
  wire [31:0] R11610;
  wire [31:0] R11609;
  wire [31:0] R11608;
  wire [31:0] R11607;
  wire [31:0] R11606;
  wire [31:0] R11605;
  wire [31:0] R11604;
  wire [31:0] R11603;
  wire [31:0] R11602;
  wire [31:0] R11601;
  wire [31:0] R11600;
  wire [31:0] R11599;
  wire [31:0] R11598;
  wire [31:0] R11597;
  wire [63:0] R11596;
  wire [31:0] R11595;
  wire [63:0] R11594;
  wire [63:0] R11593;
  wire [63:0] R11592;
  wire [63:0] R11591;
  wire [63:0] R11590;
  wire [63:0] R11589;
  wire [63:0] R11588;
  wire [63:0] R11587;
  wire [63:0] R11586;
  wire [63:0] R11585;
  wire [63:0] R11584;
  wire [63:0] R11583;
  wire [63:0] R11582;
  wire [63:0] R11581;
  wire [63:0] R11580;
  wire [63:0] R11579;
  wire [63:0] R11578;
  wire [63:0] R11577;
  wire [63:0] R11576;
  wire [63:0] R11575;
  wire [63:0] R11574;
  wire [63:0] R11573;
  wire [63:0] R11572;
  wire [63:0] R11571;
  wire [63:0] R11570;
  wire [63:0] R11569;
  wire [63:0] R11568;
  wire [63:0] R11567;
  wire [63:0] R11566;
  wire [63:0] R11565;
  wire [63:0] R11564;
  wire [63:0] R11563;
  wire [63:0] R11562;
  wire [63:0] R11561;
  wire [63:0] R11560;
  wire [63:0] R11559;
  wire [63:0] R11558;
  wire [63:0] R11557;
  wire [63:0] R11556;
  wire [63:0] R11555;
  wire [63:0] R11554;
  wire [63:0] R11553;
  wire [63:0] R11552;
  wire [63:0] R11551;
  wire [63:0] R11550;
  wire [63:0] R11549;
  wire [0:0] R11548;
  wire [0:0] R11547;
  wire [0:0] R11546;
  wire [0:0] R11545;
  wire [0:0] R11544;
  wire [0:0] R11543;
  wire [0:0] R11542;
  wire [0:0] R11541;
  wire [0:0] R11540;
  wire [0:0] R11539;
  wire [0:0] R11538;
  wire [0:0] R11537;
  wire [0:0] R11536;
  wire [0:0] R11535;
  wire [0:0] R11534;
  wire [0:0] R11533;
  wire [0:0] R11532;
  wire [0:0] R11531;
  wire [0:0] R11530;
  wire [0:0] R11529;
  wire [0:0] R11528;
  wire [0:0] R11527;
  wire [0:0] R11526;
  wire [0:0] R11525;
  wire [0:0] R11524;
  wire [0:0] R11523;
  wire [0:0] R11522;
  wire [0:0] R11521;
  wire [0:0] R11520;
  wire [0:0] R11519;
  wire [0:0] R11518;
  wire [0:0] R11517;
  wire [0:0] R11516;
  wire [0:0] R11515;
  wire [0:0] R11514;
  wire [0:0] R11513;
  wire [0:0] R11512;
  wire [0:0] R11511;
  wire [0:0] R11510;
  wire [0:0] R11509;
  wire [0:0] R11508;
  wire [0:0] R11507;
  wire [0:0] R11506;
  wire [0:0] R11505;
  wire [0:0] R11504;
  wire [0:0] R11503;
  wire [0:0] R11502;
  wire [0:0] R11501;
  wire [0:0] R11500;
  wire [0:0] R11499;
  wire [0:0] R11498;
  wire [0:0] R11497;
  wire [0:0] R11496;
  wire [0:0] R11495;
  wire [0:0] R11494;
  wire [0:0] R11493;
  wire [0:0] R11492;
  wire [0:0] R11491;
  wire [0:0] R11490;
  wire [0:0] R11489;
  wire [0:0] R11488;
  wire [0:0] R11487;
  wire [0:0] R11486;
  wire [0:0] R11485;
  wire [0:0] R11484;
  wire [0:0] R11483;
  wire [0:0] R11482;
  wire [0:0] R11481;
  wire [0:0] R11480;
  wire [0:0] R11479;
  wire [0:0] R11478;
  wire [0:0] R11477;
  wire [0:0] R11476;
  wire [0:0] R11475;
  wire [0:0] R11474;
  wire [0:0] R11473;
  wire [63:0] R11472;
  wire [31:0] R11471;
  wire [31:0] R11470;
  wire [31:0] R11469;
  wire [31:0] R11468;
  wire [31:0] R11467;
  wire [31:0] R11466;
  wire [31:0] R11465;
  wire [31:0] R11464;
  wire [31:0] R11463;
  wire [31:0] R11462;
  wire [31:0] R11461;
  wire [31:0] R11460;
  wire [31:0] R11459;
  wire [31:0] R11458;
  wire [31:0] R11457;
  wire [31:0] R11456;
  wire [31:0] R11455;
  wire [31:0] R11454;
  wire [31:0] R11453;
  wire [31:0] R11452;
  wire [31:0] R11451;
  wire [31:0] R11450;
  wire [31:0] R11449;
  wire [31:0] R11448;
  wire [31:0] R11447;
  wire [31:0] R11446;
  wire [31:0] R11445;
  wire [31:0] R11444;
  wire [31:0] R11443;
  wire [31:0] R11442;
  wire [31:0] R11441;
  wire [31:0] R11440;
  wire [31:0] R11439;
  wire [31:0] R11438;
  wire [31:0] R11437;
  wire [31:0] R11436;
  wire [31:0] R11435;
  wire [31:0] R11434;
  wire [31:0] R11433;
  wire [31:0] R11432;
  wire [31:0] R11431;
  wire [31:0] R11430;
  wire [31:0] R11429;
  wire [31:0] R11428;
  wire [31:0] R11427;
  wire [31:0] R11426;
  wire [31:0] R11425;
  wire [31:0] R11424;
  wire [31:0] R11423;
  wire [31:0] R11422;
  wire [31:0] R11421;
  wire [31:0] R11420;
  wire [31:0] R11419;
  wire [31:0] R11418;
  wire [31:0] R11417;
  wire [31:0] R11416;
  wire [31:0] R11415;
  wire [31:0] R11414;
  wire [31:0] R11413;
  wire [31:0] R11412;
  wire [31:0] R11411;
  wire [31:0] R11410;
  wire [31:0] R11409;
  wire [31:0] R11408;
  wire [31:0] R11407;
  wire [31:0] R11406;
  wire [31:0] R11405;
  wire [31:0] R11404;
  wire [31:0] R11403;
  wire [63:0] R11402;
  wire [63:0] R11401;
  wire [63:0] R11400;
  wire [31:0] R11399;
  wire [31:0] R11398;
  wire [31:0] R11397;
  wire [31:0] R11396;
  wire [31:0] R11395;
  wire [31:0] R11394;
  wire [31:0] R11393;
  wire [31:0] R11392;
  wire [31:0] R11391;
  wire [31:0] R11390;
  wire [31:0] R11389;
  wire [31:0] R11388;
  wire [31:0] R11387;
  wire [31:0] R11386;
  wire [31:0] R11385;
  wire [31:0] R11384;
  wire [31:0] R11383;
  wire [31:0] R11382;
  wire [31:0] R11381;
  wire [31:0] R11380;
  wire [31:0] R11379;
  wire [31:0] R11378;
  wire [31:0] R11377;
  wire [31:0] R11376;
  wire [31:0] R11375;
  wire [31:0] R11374;
  wire [31:0] R11373;
  wire [31:0] R11372;
  wire [31:0] R11371;
  wire [31:0] R11370;
  wire [31:0] R11369;
  wire [31:0] R11368;
  wire [31:0] R11367;
  wire [31:0] R11366;
  wire [31:0] R11365;
  wire [31:0] R11364;
  wire [31:0] R11363;
  wire [31:0] R11362;
  wire [31:0] R11361;
  wire [31:0] R11360;
  wire [31:0] R11359;
  wire [31:0] R11358;
  wire [31:0] R11357;
  wire [31:0] R11356;
  wire [31:0] R11355;
  wire [31:0] R11354;
  wire [31:0] R11353;
  wire [31:0] R11352;
  wire [31:0] R11351;
  wire [31:0] R11350;
  wire [31:0] R11349;
  wire [31:0] R11348;
  wire [31:0] R11347;
  wire [31:0] R11346;
  wire [31:0] R11345;
  wire [31:0] R11344;
  wire [31:0] R11343;
  wire [31:0] R11342;
  wire [31:0] R11341;
  wire [31:0] R11340;
  wire [31:0] R11339;
  wire [31:0] R11338;
  wire [31:0] R11337;
  wire [31:0] R11336;
  wire [31:0] R11335;
  wire [31:0] R11334;
  wire [31:0] R11333;
  wire [31:0] R11332;
  wire [31:0] R11331;
  wire [31:0] R11330;
  wire [31:0] R11329;
  wire [31:0] R11328;
  wire [31:0] R11327;
  wire [31:0] R11326;
  wire [31:0] R11325;
  wire [63:0] R11324;
  wire [31:0] R11323;
  wire [63:0] R11322;
  wire [63:0] R11321;
  wire [63:0] R11320;
  wire [63:0] R11319;
  wire [63:0] R11318;
  wire [63:0] R11317;
  wire [63:0] R11316;
  wire [63:0] R11315;
  wire [63:0] R11314;
  wire [63:0] R11313;
  wire [63:0] R11312;
  wire [63:0] R11311;
  wire [63:0] R11310;
  wire [63:0] R11309;
  wire [63:0] R11308;
  wire [63:0] R11307;
  wire [63:0] R11306;
  wire [63:0] R11305;
  wire [63:0] R11304;
  wire [63:0] R11303;
  wire [63:0] R11302;
  wire [63:0] R11301;
  wire [63:0] R11300;
  wire [63:0] R11299;
  wire [63:0] R11298;
  wire [63:0] R11297;
  wire [63:0] R11296;
  wire [63:0] R11295;
  wire [63:0] R11294;
  wire [63:0] R11293;
  wire [63:0] R11292;
  wire [63:0] R11291;
  wire [63:0] R11290;
  wire [63:0] R11289;
  wire [63:0] R11288;
  wire [63:0] R11287;
  wire [63:0] R11286;
  wire [63:0] R11285;
  wire [63:0] R11284;
  wire [63:0] R11283;
  wire [63:0] R11282;
  wire [63:0] R11281;
  wire [63:0] R11280;
  wire [63:0] R11279;
  wire [63:0] R11278;
  wire [63:0] R11277;
  wire [0:0] R11276;
  wire [0:0] R11275;
  wire [0:0] R11274;
  wire [0:0] R11273;
  wire [0:0] R11272;
  wire [0:0] R11271;
  wire [0:0] R11270;
  wire [0:0] R11269;
  wire [0:0] R11268;
  wire [0:0] R11267;
  wire [0:0] R11266;
  wire [0:0] R11265;
  wire [0:0] R11264;
  wire [0:0] R11263;
  wire [0:0] R11262;
  wire [0:0] R11261;
  wire [0:0] R11260;
  wire [0:0] R11259;
  wire [0:0] R11258;
  wire [0:0] R11257;
  wire [0:0] R11256;
  wire [0:0] R11255;
  wire [0:0] R11254;
  wire [0:0] R11253;
  wire [0:0] R11252;
  wire [0:0] R11251;
  wire [0:0] R11250;
  wire [0:0] R11249;
  wire [0:0] R11248;
  wire [0:0] R11247;
  wire [0:0] R11246;
  wire [0:0] R11245;
  wire [0:0] R11244;
  wire [0:0] R11243;
  wire [0:0] R11242;
  wire [0:0] R11241;
  wire [0:0] R11240;
  wire [0:0] R11239;
  wire [0:0] R11238;
  wire [0:0] R11237;
  wire [0:0] R11236;
  wire [0:0] R11235;
  wire [0:0] R11234;
  wire [0:0] R11233;
  wire [0:0] R11232;
  wire [0:0] R11231;
  wire [0:0] R11230;
  wire [0:0] R11229;
  wire [0:0] R11228;
  wire [0:0] R11227;
  wire [0:0] R11226;
  wire [0:0] R11225;
  wire [0:0] R11224;
  wire [0:0] R11223;
  wire [0:0] R11222;
  wire [0:0] R11221;
  wire [0:0] R11220;
  wire [0:0] R11219;
  wire [0:0] R11218;
  wire [0:0] R11217;
  wire [0:0] R11216;
  wire [0:0] R11215;
  wire [0:0] R11214;
  wire [0:0] R11213;
  wire [0:0] R11212;
  wire [0:0] R11211;
  wire [0:0] R11210;
  wire [0:0] R11209;
  wire [0:0] R11208;
  wire [0:0] R11207;
  wire [0:0] R11206;
  wire [0:0] R11205;
  wire [0:0] R11204;
  wire [0:0] R11203;
  wire [0:0] R11202;
  wire [0:0] R11201;
  wire [0:0] R11200;
  wire [0:0] R11199;
  wire [0:0] R11198;
  wire [0:0] R11197;
  wire [0:0] R11196;
  wire [0:0] R11195;
  wire [0:0] R11194;
  wire [0:0] R11193;
  wire [0:0] R11192;
  wire [0:0] R11191;
  wire [0:0] R11190;
  wire [0:0] R11189;
  wire [0:0] R11188;
  wire [63:0] R11187;
  wire [31:0] R11186;
  wire [31:0] R11185;
  wire [31:0] R11184;
  wire [31:0] R11183;
  wire [31:0] R11182;
  wire [31:0] R11181;
  wire [31:0] R11180;
  wire [31:0] R11179;
  wire [31:0] R11178;
  wire [31:0] R11177;
  wire [31:0] R11176;
  wire [31:0] R11175;
  wire [31:0] R11174;
  wire [31:0] R11173;
  wire [31:0] R11172;
  wire [31:0] R11171;
  wire [31:0] R11170;
  wire [31:0] R11169;
  wire [31:0] R11168;
  wire [31:0] R11167;
  wire [31:0] R11166;
  wire [31:0] R11165;
  wire [31:0] R11164;
  wire [31:0] R11163;
  wire [31:0] R11162;
  wire [31:0] R11161;
  wire [31:0] R11160;
  wire [31:0] R11159;
  wire [31:0] R11158;
  wire [31:0] R11157;
  wire [31:0] R11156;
  wire [31:0] R11155;
  wire [31:0] R11154;
  wire [31:0] R11153;
  wire [31:0] R11152;
  wire [31:0] R11151;
  wire [31:0] R11150;
  wire [31:0] R11149;
  wire [31:0] R11148;
  wire [31:0] R11147;
  wire [31:0] R11146;
  wire [31:0] R11145;
  wire [31:0] R11144;
  wire [31:0] R11143;
  wire [31:0] R11142;
  wire [31:0] R11141;
  wire [31:0] R11140;
  wire [31:0] R11139;
  wire [31:0] R11138;
  wire [31:0] R11137;
  wire [31:0] R11136;
  wire [31:0] R11135;
  wire [31:0] R11134;
  wire [31:0] R11133;
  wire [31:0] R11132;
  wire [31:0] R11131;
  wire [31:0] R11130;
  wire [31:0] R11129;
  wire [31:0] R11128;
  wire [31:0] R11127;
  wire [31:0] R11126;
  wire [31:0] R11125;
  wire [31:0] R11124;
  wire [31:0] R11123;
  wire [31:0] R11122;
  wire [31:0] R11121;
  wire [31:0] R11120;
  wire [31:0] R11119;
  wire [31:0] R11118;
  wire [31:0] R11117;
  wire [31:0] R11116;
  wire [31:0] R11115;
  wire [31:0] R11114;
  wire [31:0] R11113;
  wire [31:0] R11112;
  wire [31:0] R11111;
  wire [31:0] R11110;
  wire [31:0] R11109;
  wire [31:0] R11108;
  wire [31:0] R11107;
  wire [31:0] R11106;
  wire [31:0] R11105;
  wire [63:0] R11104;
  wire [63:0] R11103;
  wire [63:0] R11102;
  wire [31:0] R11101;
  wire [31:0] R11100;
  wire [31:0] R11099;
  wire [31:0] R11098;
  wire [31:0] R11097;
  wire [31:0] R11096;
  wire [31:0] R11095;
  wire [31:0] R11094;
  wire [31:0] R11093;
  wire [31:0] R11092;
  wire [31:0] R11091;
  wire [31:0] R11090;
  wire [31:0] R11089;
  wire [31:0] R11088;
  wire [31:0] R11087;
  wire [31:0] R11086;
  wire [31:0] R11085;
  wire [31:0] R11084;
  wire [31:0] R11083;
  wire [31:0] R11082;
  wire [31:0] R11081;
  wire [31:0] R11080;
  wire [31:0] R11079;
  wire [31:0] R11078;
  wire [31:0] R11077;
  wire [31:0] R11076;
  wire [31:0] R11075;
  wire [31:0] R11074;
  wire [31:0] R11073;
  wire [31:0] R11072;
  wire [31:0] R11071;
  wire [31:0] R11070;
  wire [31:0] R11069;
  wire [31:0] R11068;
  wire [31:0] R11067;
  wire [31:0] R11066;
  wire [31:0] R11065;
  wire [31:0] R11064;
  wire [31:0] R11063;
  wire [31:0] R11062;
  wire [31:0] R11061;
  wire [31:0] R11060;
  wire [31:0] R11059;
  wire [31:0] R11058;
  wire [31:0] R11057;
  wire [31:0] R11056;
  wire [31:0] R11055;
  wire [31:0] R11054;
  wire [31:0] R11053;
  wire [31:0] R11052;
  wire [31:0] R11051;
  wire [31:0] R11050;
  wire [31:0] R11049;
  wire [31:0] R11048;
  wire [31:0] R11047;
  wire [31:0] R11046;
  wire [31:0] R11045;
  wire [31:0] R11044;
  wire [31:0] R11043;
  wire [31:0] R11042;
  wire [31:0] R11041;
  wire [31:0] R11040;
  wire [31:0] R11039;
  wire [31:0] R11038;
  wire [31:0] R11037;
  wire [31:0] R11036;
  wire [31:0] R11035;
  wire [31:0] R11034;
  wire [31:0] R11033;
  wire [31:0] R11032;
  wire [31:0] R11031;
  wire [31:0] R11030;
  wire [31:0] R11029;
  wire [31:0] R11028;
  wire [31:0] R11027;
  wire [31:0] R11026;
  wire [31:0] R11025;
  wire [31:0] R11024;
  wire [31:0] R11023;
  wire [31:0] R11022;
  wire [31:0] R11021;
  wire [31:0] R11020;
  wire [31:0] R11019;
  wire [31:0] R11018;
  wire [31:0] R11017;
  wire [31:0] R11016;
  wire [31:0] R11015;
  wire [31:0] R11014;
  wire [63:0] R11013;
  wire [31:0] R11012;
  wire [63:0] R11011;
  wire [63:0] R11010;
  wire [63:0] R11009;
  wire [63:0] R11008;
  wire [63:0] R11007;
  wire [63:0] R11006;
  wire [63:0] R11005;
  wire [63:0] R11004;
  wire [63:0] R11003;
  wire [63:0] R11002;
  wire [63:0] R11001;
  wire [63:0] R11000;
  wire [63:0] R10999;
  wire [63:0] R10998;
  wire [63:0] R10997;
  wire [63:0] R10996;
  wire [63:0] R10995;
  wire [63:0] R10994;
  wire [63:0] R10993;
  wire [63:0] R10992;
  wire [63:0] R10991;
  wire [63:0] R10990;
  wire [63:0] R10989;
  wire [63:0] R10988;
  wire [63:0] R10987;
  wire [63:0] R10986;
  wire [63:0] R10985;
  wire [63:0] R10984;
  wire [63:0] R10983;
  wire [63:0] R10982;
  wire [63:0] R10981;
  wire [63:0] R10980;
  wire [63:0] R10979;
  wire [63:0] R10978;
  wire [63:0] R10977;
  wire [63:0] R10976;
  wire [63:0] R10975;
  wire [63:0] R10974;
  wire [63:0] R10973;
  wire [63:0] R10972;
  wire [63:0] R10971;
  wire [63:0] R10970;
  wire [63:0] R10969;
  wire [63:0] R10968;
  wire [63:0] R10967;
  wire [63:0] R10966;
  wire [0:0] R10965;
  wire [0:0] R10964;
  wire [0:0] R10963;
  wire [0:0] R10962;
  wire [0:0] R10961;
  wire [0:0] R10960;
  wire [0:0] R10959;
  wire [0:0] R10958;
  wire [0:0] R10957;
  wire [0:0] R10956;
  wire [0:0] R10955;
  wire [0:0] R10954;
  wire [0:0] R10953;
  wire [0:0] R10952;
  wire [0:0] R10951;
  wire [0:0] R10950;
  wire [0:0] R10949;
  wire [0:0] R10948;
  wire [0:0] R10947;
  wire [0:0] R10946;
  wire [0:0] R10945;
  wire [0:0] R10944;
  wire [0:0] R10943;
  wire [0:0] R10942;
  wire [0:0] R10941;
  wire [0:0] R10940;
  wire [0:0] R10939;
  wire [0:0] R10938;
  wire [0:0] R10937;
  wire [0:0] R10936;
  wire [0:0] R10935;
  wire [0:0] R10934;
  wire [0:0] R10933;
  wire [0:0] R10932;
  wire [0:0] R10931;
  wire [0:0] R10930;
  wire [0:0] R10929;
  wire [0:0] R10928;
  wire [0:0] R10927;
  wire [0:0] R10926;
  wire [0:0] R10925;
  wire [0:0] R10924;
  wire [0:0] R10923;
  wire [0:0] R10922;
  wire [0:0] R10921;
  wire [0:0] R10920;
  wire [0:0] R10919;
  wire [0:0] R10918;
  wire [0:0] R10917;
  wire [0:0] R10916;
  wire [0:0] R10915;
  wire [0:0] R10914;
  wire [0:0] R10913;
  wire [0:0] R10912;
  wire [0:0] R10911;
  wire [0:0] R10910;
  wire [0:0] R10909;
  wire [0:0] R10908;
  wire [0:0] R10907;
  wire [0:0] R10906;
  wire [0:0] R10905;
  wire [0:0] R10904;
  wire [0:0] R10903;
  wire [0:0] R10902;
  wire [0:0] R10901;
  wire [0:0] R10900;
  wire [0:0] R10899;
  wire [0:0] R10898;
  wire [0:0] R10897;
  wire [0:0] R10896;
  wire [0:0] R10895;
  wire [0:0] R10894;
  wire [0:0] R10893;
  wire [0:0] R10892;
  wire [0:0] R10891;
  wire [0:0] R10890;
  wire [0:0] R10889;
  wire [0:0] R10888;
  wire [0:0] R10887;
  wire [0:0] R10886;
  wire [0:0] R10885;
  wire [0:0] R10884;
  wire [0:0] R10883;
  wire [0:0] R10882;
  wire [0:0] R10881;
  wire [0:0] R10880;
  wire [0:0] R10879;
  wire [0:0] R10878;
  wire [0:0] R10877;
  wire [0:0] R10876;
  wire [0:0] R10875;
  wire [0:0] R10874;
  wire [0:0] R10873;
  wire [0:0] R10872;
  wire [0:0] R10871;
  wire [0:0] R10870;
  wire [0:0] R10869;
  wire [0:0] R10868;
  wire [0:0] R10867;
  wire [0:0] R10866;
  wire [0:0] R10865;
  wire [0:0] R10864;
  wire [63:0] R10863;
  wire [31:0] R10862;
  wire [31:0] R10861;
  wire [31:0] R10860;
  wire [31:0] R10859;
  wire [31:0] R10858;
  wire [31:0] R10857;
  wire [31:0] R10856;
  wire [31:0] R10855;
  wire [31:0] R10854;
  wire [31:0] R10853;
  wire [31:0] R10852;
  wire [31:0] R10851;
  wire [31:0] R10850;
  wire [31:0] R10849;
  wire [31:0] R10848;
  wire [31:0] R10847;
  wire [31:0] R10846;
  wire [31:0] R10845;
  wire [31:0] R10844;
  wire [31:0] R10843;
  wire [31:0] R10842;
  wire [31:0] R10841;
  wire [31:0] R10840;
  wire [31:0] R10839;
  wire [31:0] R10838;
  wire [31:0] R10837;
  wire [31:0] R10836;
  wire [31:0] R10835;
  wire [31:0] R10834;
  wire [31:0] R10833;
  wire [31:0] R10832;
  wire [31:0] R10831;
  wire [31:0] R10830;
  wire [31:0] R10829;
  wire [31:0] R10828;
  wire [31:0] R10827;
  wire [31:0] R10826;
  wire [31:0] R10825;
  wire [31:0] R10824;
  wire [31:0] R10823;
  wire [31:0] R10822;
  wire [31:0] R10821;
  wire [31:0] R10820;
  wire [31:0] R10819;
  wire [31:0] R10818;
  wire [31:0] R10817;
  wire [31:0] R10816;
  wire [31:0] R10815;
  wire [31:0] R10814;
  wire [31:0] R10813;
  wire [31:0] R10812;
  wire [31:0] R10811;
  wire [31:0] R10810;
  wire [31:0] R10809;
  wire [31:0] R10808;
  wire [31:0] R10807;
  wire [31:0] R10806;
  wire [31:0] R10805;
  wire [31:0] R10804;
  wire [31:0] R10803;
  wire [31:0] R10802;
  wire [31:0] R10801;
  wire [31:0] R10800;
  wire [31:0] R10799;
  wire [31:0] R10798;
  wire [31:0] R10797;
  wire [31:0] R10796;
  wire [31:0] R10795;
  wire [31:0] R10794;
  wire [31:0] R10793;
  wire [31:0] R10792;
  wire [31:0] R10791;
  wire [31:0] R10790;
  wire [31:0] R10789;
  wire [31:0] R10788;
  wire [31:0] R10787;
  wire [31:0] R10786;
  wire [31:0] R10785;
  wire [31:0] R10784;
  wire [31:0] R10783;
  wire [31:0] R10782;
  wire [31:0] R10781;
  wire [31:0] R10780;
  wire [31:0] R10779;
  wire [31:0] R10778;
  wire [31:0] R10777;
  wire [31:0] R10776;
  wire [31:0] R10775;
  wire [31:0] R10774;
  wire [31:0] R10773;
  wire [31:0] R10772;
  wire [31:0] R10771;
  wire [31:0] R10770;
  wire [31:0] R10769;
  wire [31:0] R10768;
  wire [63:0] R10767;
  wire [63:0] R10766;
  wire [63:0] R10765;
  wire [31:0] R10764;
  wire [31:0] R10763;
  wire [31:0] R10762;
  wire [31:0] R10761;
  wire [31:0] R10760;
  wire [31:0] R10759;
  wire [31:0] R10758;
  wire [31:0] R10757;
  wire [31:0] R10756;
  wire [31:0] R10755;
  wire [31:0] R10754;
  wire [31:0] R10753;
  wire [31:0] R10752;
  wire [31:0] R10751;
  wire [31:0] R10750;
  wire [31:0] R10749;
  wire [31:0] R10748;
  wire [31:0] R10747;
  wire [31:0] R10746;
  wire [31:0] R10745;
  wire [31:0] R10744;
  wire [31:0] R10743;
  wire [31:0] R10742;
  wire [31:0] R10741;
  wire [31:0] R10740;
  wire [31:0] R10739;
  wire [31:0] R10738;
  wire [31:0] R10737;
  wire [31:0] R10736;
  wire [31:0] R10735;
  wire [31:0] R10734;
  wire [31:0] R10733;
  wire [31:0] R10732;
  wire [31:0] R10731;
  wire [31:0] R10730;
  wire [31:0] R10729;
  wire [31:0] R10728;
  wire [31:0] R10727;
  wire [31:0] R10726;
  wire [31:0] R10725;
  wire [31:0] R10724;
  wire [31:0] R10723;
  wire [31:0] R10722;
  wire [31:0] R10721;
  wire [31:0] R10720;
  wire [31:0] R10719;
  wire [31:0] R10718;
  wire [31:0] R10717;
  wire [31:0] R10716;
  wire [31:0] R10715;
  wire [31:0] R10714;
  wire [31:0] R10713;
  wire [31:0] R10712;
  wire [31:0] R10711;
  wire [31:0] R10710;
  wire [31:0] R10709;
  wire [31:0] R10708;
  wire [31:0] R10707;
  wire [31:0] R10706;
  wire [31:0] R10705;
  wire [31:0] R10704;
  wire [31:0] R10703;
  wire [31:0] R10702;
  wire [31:0] R10701;
  wire [31:0] R10700;
  wire [31:0] R10699;
  wire [31:0] R10698;
  wire [31:0] R10697;
  wire [31:0] R10696;
  wire [31:0] R10695;
  wire [31:0] R10694;
  wire [31:0] R10693;
  wire [31:0] R10692;
  wire [31:0] R10691;
  wire [31:0] R10690;
  wire [31:0] R10689;
  wire [31:0] R10688;
  wire [31:0] R10687;
  wire [31:0] R10686;
  wire [31:0] R10685;
  wire [31:0] R10684;
  wire [31:0] R10683;
  wire [31:0] R10682;
  wire [31:0] R10681;
  wire [31:0] R10680;
  wire [31:0] R10679;
  wire [31:0] R10678;
  wire [31:0] R10677;
  wire [31:0] R10676;
  wire [31:0] R10675;
  wire [31:0] R10674;
  wire [31:0] R10673;
  wire [31:0] R10672;
  wire [31:0] R10671;
  wire [31:0] R10670;
  wire [31:0] R10669;
  wire [31:0] R10668;
  wire [31:0] R10667;
  wire [31:0] R10666;
  wire [31:0] R10665;
  wire [31:0] R10664;
  wire [63:0] R10663;
  wire [31:0] R10662;
  wire [63:0] R10661;
  wire [63:0] R10660;
  wire [63:0] R10659;
  wire [63:0] R10658;
  wire [63:0] R10657;
  wire [63:0] R10656;
  wire [63:0] R10655;
  wire [63:0] R10654;
  wire [63:0] R10653;
  wire [63:0] R10652;
  wire [63:0] R10651;
  wire [63:0] R10650;
  wire [63:0] R10649;
  wire [63:0] R10648;
  wire [63:0] R10647;
  wire [63:0] R10646;
  wire [63:0] R10645;
  wire [63:0] R10644;
  wire [63:0] R10643;
  wire [63:0] R10642;
  wire [63:0] R10641;
  wire [63:0] R10640;
  wire [63:0] R10639;
  wire [63:0] R10638;
  wire [63:0] R10637;
  wire [63:0] R10636;
  wire [63:0] R10635;
  wire [63:0] R10634;
  wire [63:0] R10633;
  wire [63:0] R10632;
  wire [63:0] R10631;
  wire [63:0] R10630;
  wire [63:0] R10629;
  wire [63:0] R10628;
  wire [63:0] R10627;
  wire [63:0] R10626;
  wire [63:0] R10625;
  wire [63:0] R10624;
  wire [63:0] R10623;
  wire [63:0] R10622;
  wire [63:0] R10621;
  wire [63:0] R10620;
  wire [63:0] R10619;
  wire [63:0] R10618;
  wire [63:0] R10617;
  wire [63:0] R10616;
  wire [0:0] R10615;
  wire [0:0] R10614;
  wire [0:0] R10613;
  wire [0:0] R10612;
  wire [0:0] R10611;
  wire [0:0] R10610;
  wire [0:0] R10609;
  wire [0:0] R10608;
  wire [0:0] R10607;
  wire [0:0] R10606;
  wire [0:0] R10605;
  wire [0:0] R10604;
  wire [0:0] R10603;
  wire [0:0] R10602;
  wire [0:0] R10601;
  wire [0:0] R10600;
  wire [0:0] R10599;
  wire [0:0] R10598;
  wire [0:0] R10597;
  wire [0:0] R10596;
  wire [0:0] R10595;
  wire [0:0] R10594;
  wire [0:0] R10593;
  wire [0:0] R10592;
  wire [0:0] R10591;
  wire [0:0] R10590;
  wire [0:0] R10589;
  wire [0:0] R10588;
  wire [0:0] R10587;
  wire [0:0] R10586;
  wire [0:0] R10585;
  wire [0:0] R10584;
  wire [0:0] R10583;
  wire [0:0] R10582;
  wire [0:0] R10581;
  wire [0:0] R10580;
  wire [0:0] R10579;
  wire [0:0] R10578;
  wire [0:0] R10577;
  wire [0:0] R10576;
  wire [0:0] R10575;
  wire [0:0] R10574;
  wire [0:0] R10573;
  wire [0:0] R10572;
  wire [0:0] R10571;
  wire [0:0] R10570;
  wire [0:0] R10569;
  wire [0:0] R10568;
  wire [0:0] R10567;
  wire [0:0] R10566;
  wire [0:0] R10565;
  wire [0:0] R10564;
  wire [0:0] R10563;
  wire [0:0] R10562;
  wire [0:0] R10561;
  wire [0:0] R10560;
  wire [0:0] R10559;
  wire [0:0] R10558;
  wire [0:0] R10557;
  wire [0:0] R10556;
  wire [0:0] R10555;
  wire [0:0] R10554;
  wire [0:0] R10553;
  wire [0:0] R10552;
  wire [0:0] R10551;
  wire [0:0] R10550;
  wire [0:0] R10549;
  wire [0:0] R10548;
  wire [0:0] R10547;
  wire [0:0] R10546;
  wire [0:0] R10545;
  wire [0:0] R10544;
  wire [0:0] R10543;
  wire [0:0] R10542;
  wire [0:0] R10541;
  wire [0:0] R10540;
  wire [0:0] R10539;
  wire [0:0] R10538;
  wire [0:0] R10537;
  wire [0:0] R10536;
  wire [0:0] R10535;
  wire [0:0] R10534;
  wire [0:0] R10533;
  wire [0:0] R10532;
  wire [0:0] R10531;
  wire [0:0] R10530;
  wire [0:0] R10529;
  wire [0:0] R10528;
  wire [0:0] R10527;
  wire [0:0] R10526;
  wire [0:0] R10525;
  wire [0:0] R10524;
  wire [0:0] R10523;
  wire [0:0] R10522;
  wire [0:0] R10521;
  wire [0:0] R10520;
  wire [0:0] R10519;
  wire [0:0] R10518;
  wire [0:0] R10517;
  wire [0:0] R10516;
  wire [0:0] R10515;
  wire [0:0] R10514;
  wire [0:0] R10513;
  wire [0:0] R10512;
  wire [0:0] R10511;
  wire [0:0] R10510;
  wire [0:0] R10509;
  wire [0:0] R10508;
  wire [0:0] R10507;
  wire [0:0] R10506;
  wire [0:0] R10505;
  wire [0:0] R10504;
  wire [0:0] R10503;
  wire [0:0] R10502;
  wire [0:0] R10501;
  wire [0:0] R10500;
  wire [63:0] R10499;
  wire [31:0] R10498;
  wire [31:0] R10497;
  wire [31:0] R10496;
  wire [31:0] R10495;
  wire [31:0] R10494;
  wire [31:0] R10493;
  wire [31:0] R10492;
  wire [31:0] R10491;
  wire [31:0] R10490;
  wire [31:0] R10489;
  wire [31:0] R10488;
  wire [31:0] R10487;
  wire [31:0] R10486;
  wire [31:0] R10485;
  wire [31:0] R10484;
  wire [31:0] R10483;
  wire [31:0] R10482;
  wire [31:0] R10481;
  wire [31:0] R10480;
  wire [31:0] R10479;
  wire [31:0] R10478;
  wire [31:0] R10477;
  wire [31:0] R10476;
  wire [31:0] R10475;
  wire [31:0] R10474;
  wire [31:0] R10473;
  wire [31:0] R10472;
  wire [31:0] R10471;
  wire [31:0] R10470;
  wire [31:0] R10469;
  wire [31:0] R10468;
  wire [31:0] R10467;
  wire [31:0] R10466;
  wire [31:0] R10465;
  wire [31:0] R10464;
  wire [31:0] R10463;
  wire [31:0] R10462;
  wire [31:0] R10461;
  wire [31:0] R10460;
  wire [31:0] R10459;
  wire [31:0] R10458;
  wire [31:0] R10457;
  wire [31:0] R10456;
  wire [31:0] R10455;
  wire [31:0] R10454;
  wire [31:0] R10453;
  wire [31:0] R10452;
  wire [31:0] R10451;
  wire [31:0] R10450;
  wire [31:0] R10449;
  wire [31:0] R10448;
  wire [31:0] R10447;
  wire [31:0] R10446;
  wire [31:0] R10445;
  wire [31:0] R10444;
  wire [31:0] R10443;
  wire [31:0] R10442;
  wire [31:0] R10441;
  wire [31:0] R10440;
  wire [31:0] R10439;
  wire [31:0] R10438;
  wire [31:0] R10437;
  wire [31:0] R10436;
  wire [31:0] R10435;
  wire [31:0] R10434;
  wire [31:0] R10433;
  wire [31:0] R10432;
  wire [31:0] R10431;
  wire [31:0] R10430;
  wire [31:0] R10429;
  wire [31:0] R10428;
  wire [31:0] R10427;
  wire [31:0] R10426;
  wire [31:0] R10425;
  wire [31:0] R10424;
  wire [31:0] R10423;
  wire [31:0] R10422;
  wire [31:0] R10421;
  wire [31:0] R10420;
  wire [31:0] R10419;
  wire [31:0] R10418;
  wire [31:0] R10417;
  wire [31:0] R10416;
  wire [31:0] R10415;
  wire [31:0] R10414;
  wire [31:0] R10413;
  wire [31:0] R10412;
  wire [31:0] R10411;
  wire [31:0] R10410;
  wire [31:0] R10409;
  wire [31:0] R10408;
  wire [31:0] R10407;
  wire [31:0] R10406;
  wire [31:0] R10405;
  wire [31:0] R10404;
  wire [31:0] R10403;
  wire [31:0] R10402;
  wire [31:0] R10401;
  wire [31:0] R10400;
  wire [31:0] R10399;
  wire [31:0] R10398;
  wire [31:0] R10397;
  wire [31:0] R10396;
  wire [31:0] R10395;
  wire [31:0] R10394;
  wire [31:0] R10393;
  wire [31:0] R10392;
  wire [31:0] R10391;
  wire [63:0] R10390;
  wire [63:0] R10389;
  wire [63:0] R10388;
  wire [31:0] R10387;
  wire [31:0] R10386;
  wire [31:0] R10385;
  wire [31:0] R10384;
  wire [31:0] R10383;
  wire [31:0] R10382;
  wire [31:0] R10381;
  wire [31:0] R10380;
  wire [31:0] R10379;
  wire [31:0] R10378;
  wire [31:0] R10377;
  wire [31:0] R10376;
  wire [31:0] R10375;
  wire [31:0] R10374;
  wire [31:0] R10373;
  wire [31:0] R10372;
  wire [31:0] R10371;
  wire [31:0] R10370;
  wire [31:0] R10369;
  wire [31:0] R10368;
  wire [31:0] R10367;
  wire [31:0] R10366;
  wire [31:0] R10365;
  wire [31:0] R10364;
  wire [31:0] R10363;
  wire [31:0] R10362;
  wire [31:0] R10361;
  wire [31:0] R10360;
  wire [31:0] R10359;
  wire [31:0] R10358;
  wire [31:0] R10357;
  wire [31:0] R10356;
  wire [31:0] R10355;
  wire [31:0] R10354;
  wire [31:0] R10353;
  wire [31:0] R10352;
  wire [31:0] R10351;
  wire [31:0] R10350;
  wire [31:0] R10349;
  wire [31:0] R10348;
  wire [31:0] R10347;
  wire [31:0] R10346;
  wire [31:0] R10345;
  wire [31:0] R10344;
  wire [31:0] R10343;
  wire [31:0] R10342;
  wire [31:0] R10341;
  wire [31:0] R10340;
  wire [31:0] R10339;
  wire [31:0] R10338;
  wire [31:0] R10337;
  wire [31:0] R10336;
  wire [31:0] R10335;
  wire [31:0] R10334;
  wire [31:0] R10333;
  wire [31:0] R10332;
  wire [31:0] R10331;
  wire [31:0] R10330;
  wire [31:0] R10329;
  wire [31:0] R10328;
  wire [31:0] R10327;
  wire [31:0] R10326;
  wire [31:0] R10325;
  wire [31:0] R10324;
  wire [31:0] R10323;
  wire [31:0] R10322;
  wire [31:0] R10321;
  wire [31:0] R10320;
  wire [31:0] R10319;
  wire [31:0] R10318;
  wire [31:0] R10317;
  wire [31:0] R10316;
  wire [31:0] R10315;
  wire [31:0] R10314;
  wire [31:0] R10313;
  wire [31:0] R10312;
  wire [31:0] R10311;
  wire [31:0] R10310;
  wire [31:0] R10309;
  wire [31:0] R10308;
  wire [31:0] R10307;
  wire [31:0] R10306;
  wire [31:0] R10305;
  wire [31:0] R10304;
  wire [31:0] R10303;
  wire [31:0] R10302;
  wire [31:0] R10301;
  wire [31:0] R10300;
  wire [31:0] R10299;
  wire [31:0] R10298;
  wire [31:0] R10297;
  wire [31:0] R10296;
  wire [31:0] R10295;
  wire [31:0] R10294;
  wire [31:0] R10293;
  wire [31:0] R10292;
  wire [31:0] R10291;
  wire [31:0] R10290;
  wire [31:0] R10289;
  wire [31:0] R10288;
  wire [31:0] R10287;
  wire [31:0] R10286;
  wire [31:0] R10285;
  wire [31:0] R10284;
  wire [31:0] R10283;
  wire [31:0] R10282;
  wire [31:0] R10281;
  wire [31:0] R10280;
  wire [31:0] R10279;
  wire [31:0] R10278;
  wire [31:0] R10277;
  wire [31:0] R10276;
  wire [31:0] R10275;
  wire [31:0] R10274;
  wire [63:0] R10273;
  wire [31:0] R10272;
  wire [63:0] R10271;
  wire [63:0] R10270;
  wire [63:0] R10269;
  wire [63:0] R10268;
  wire [63:0] R10267;
  wire [63:0] R10266;
  wire [63:0] R10265;
  wire [63:0] R10264;
  wire [63:0] R10263;
  wire [63:0] R10262;
  wire [63:0] R10261;
  wire [63:0] R10260;
  wire [63:0] R10259;
  wire [63:0] R10258;
  wire [63:0] R10257;
  wire [63:0] R10256;
  wire [63:0] R10255;
  wire [63:0] R10254;
  wire [63:0] R10253;
  wire [63:0] R10252;
  wire [63:0] R10251;
  wire [63:0] R10250;
  wire [63:0] R10249;
  wire [63:0] R10248;
  wire [63:0] R10247;
  wire [63:0] R10246;
  wire [63:0] R10245;
  wire [63:0] R10244;
  wire [63:0] R10243;
  wire [63:0] R10242;
  wire [63:0] R10241;
  wire [63:0] R10240;
  wire [63:0] R10239;
  wire [63:0] R10238;
  wire [63:0] R10237;
  wire [63:0] R10236;
  wire [63:0] R10235;
  wire [63:0] R10234;
  wire [63:0] R10233;
  wire [63:0] R10232;
  wire [63:0] R10231;
  wire [63:0] R10230;
  wire [63:0] R10229;
  wire [63:0] R10228;
  wire [63:0] R10227;
  wire [63:0] R10226;
  wire [0:0] R10225;
  wire [0:0] R10224;
  wire [0:0] R10223;
  wire [0:0] R10222;
  wire [0:0] R10221;
  wire [0:0] R10220;
  wire [0:0] R10219;
  wire [0:0] R10218;
  wire [0:0] R10217;
  wire [0:0] R10216;
  wire [0:0] R10215;
  wire [0:0] R10214;
  wire [0:0] R10213;
  wire [0:0] R10212;
  wire [0:0] R10211;
  wire [0:0] R10210;
  wire [0:0] R10209;
  wire [0:0] R10208;
  wire [0:0] R10207;
  wire [0:0] R10206;
  wire [0:0] R10205;
  wire [0:0] R10204;
  wire [0:0] R10203;
  wire [0:0] R10202;
  wire [0:0] R10201;
  wire [0:0] R10200;
  wire [0:0] R10199;
  wire [0:0] R10198;
  wire [0:0] R10197;
  wire [0:0] R10196;
  wire [0:0] R10195;
  wire [0:0] R10194;
  wire [0:0] R10193;
  wire [0:0] R10192;
  wire [0:0] R10191;
  wire [0:0] R10190;
  wire [0:0] R10189;
  wire [0:0] R10188;
  wire [0:0] R10187;
  wire [0:0] R10186;
  wire [0:0] R10185;
  wire [0:0] R10184;
  wire [0:0] R10183;
  wire [0:0] R10182;
  wire [0:0] R10181;
  wire [0:0] R10180;
  wire [0:0] R10179;
  wire [0:0] R10178;
  wire [0:0] R10177;
  wire [0:0] R10176;
  wire [0:0] R10175;
  wire [0:0] R10174;
  wire [0:0] R10173;
  wire [0:0] R10172;
  wire [0:0] R10171;
  wire [0:0] R10170;
  wire [0:0] R10169;
  wire [0:0] R10168;
  wire [0:0] R10167;
  wire [0:0] R10166;
  wire [0:0] R10165;
  wire [0:0] R10164;
  wire [0:0] R10163;
  wire [0:0] R10162;
  wire [0:0] R10161;
  wire [0:0] R10160;
  wire [0:0] R10159;
  wire [0:0] R10158;
  wire [0:0] R10157;
  wire [0:0] R10156;
  wire [0:0] R10155;
  wire [0:0] R10154;
  wire [0:0] R10153;
  wire [0:0] R10152;
  wire [0:0] R10151;
  wire [0:0] R10150;
  wire [0:0] R10149;
  wire [0:0] R10148;
  wire [0:0] R10147;
  wire [0:0] R10146;
  wire [0:0] R10145;
  wire [0:0] R10144;
  wire [0:0] R10143;
  wire [0:0] R10142;
  wire [0:0] R10141;
  wire [0:0] R10140;
  wire [0:0] R10139;
  wire [0:0] R10138;
  wire [0:0] R10137;
  wire [0:0] R10136;
  wire [0:0] R10135;
  wire [0:0] R10134;
  wire [0:0] R10133;
  wire [0:0] R10132;
  wire [0:0] R10131;
  wire [0:0] R10130;
  wire [0:0] R10129;
  wire [0:0] R10128;
  wire [0:0] R10127;
  wire [0:0] R10126;
  wire [0:0] R10125;
  wire [0:0] R10124;
  wire [0:0] R10123;
  wire [0:0] R10122;
  wire [0:0] R10121;
  wire [0:0] R10120;
  wire [0:0] R10119;
  wire [0:0] R10118;
  wire [0:0] R10117;
  wire [0:0] R10116;
  wire [0:0] R10115;
  wire [0:0] R10114;
  wire [0:0] R10113;
  wire [0:0] R10112;
  wire [0:0] R10111;
  wire [0:0] R10110;
  wire [0:0] R10109;
  wire [0:0] R10108;
  wire [0:0] R10107;
  wire [0:0] R10106;
  wire [0:0] R10105;
  wire [0:0] R10104;
  wire [0:0] R10103;
  wire [0:0] R10102;
  wire [0:0] R10101;
  wire [0:0] R10100;
  wire [0:0] R10099;
  wire [0:0] R10098;
  wire [0:0] R10097;
  wire [63:0] R10096;
  wire [31:0] R10095;
  wire [31:0] R10094;
  wire [31:0] R10093;
  wire [31:0] R10092;
  wire [31:0] R10091;
  wire [31:0] R10090;
  wire [31:0] R10089;
  wire [31:0] R10088;
  wire [31:0] R10087;
  wire [31:0] R10086;
  wire [31:0] R10085;
  wire [31:0] R10084;
  wire [31:0] R10083;
  wire [31:0] R10082;
  wire [31:0] R10081;
  wire [31:0] R10080;
  wire [31:0] R10079;
  wire [31:0] R10078;
  wire [31:0] R10077;
  wire [31:0] R10076;
  wire [31:0] R10075;
  wire [31:0] R10074;
  wire [31:0] R10073;
  wire [31:0] R10072;
  wire [31:0] R10071;
  wire [31:0] R10070;
  wire [31:0] R10069;
  wire [31:0] R10068;
  wire [31:0] R10067;
  wire [31:0] R10066;
  wire [31:0] R10065;
  wire [31:0] R10064;
  wire [31:0] R10063;
  wire [31:0] R10062;
  wire [31:0] R10061;
  wire [31:0] R10060;
  wire [31:0] R10059;
  wire [31:0] R10058;
  wire [31:0] R10057;
  wire [31:0] R10056;
  wire [31:0] R10055;
  wire [31:0] R10054;
  wire [31:0] R10053;
  wire [31:0] R10052;
  wire [31:0] R10051;
  wire [31:0] R10050;
  wire [31:0] R10049;
  wire [31:0] R10048;
  wire [31:0] R10047;
  wire [31:0] R10046;
  wire [31:0] R10045;
  wire [31:0] R10044;
  wire [31:0] R10043;
  wire [31:0] R10042;
  wire [31:0] R10041;
  wire [31:0] R10040;
  wire [31:0] R10039;
  wire [31:0] R10038;
  wire [31:0] R10037;
  wire [31:0] R10036;
  wire [31:0] R10035;
  wire [31:0] R10034;
  wire [31:0] R10033;
  wire [31:0] R10032;
  wire [31:0] R10031;
  wire [31:0] R10030;
  wire [31:0] R10029;
  wire [31:0] R10028;
  wire [31:0] R10027;
  wire [31:0] R10026;
  wire [31:0] R10025;
  wire [31:0] R10024;
  wire [31:0] R10023;
  wire [31:0] R10022;
  wire [31:0] R10021;
  wire [31:0] R10020;
  wire [31:0] R10019;
  wire [31:0] R10018;
  wire [31:0] R10017;
  wire [31:0] R10016;
  wire [31:0] R10015;
  wire [31:0] R10014;
  wire [31:0] R10013;
  wire [31:0] R10012;
  wire [31:0] R10011;
  wire [31:0] R10010;
  wire [31:0] R10009;
  wire [31:0] R10008;
  wire [31:0] R10007;
  wire [31:0] R10006;
  wire [31:0] R10005;
  wire [31:0] R10004;
  wire [31:0] R10003;
  wire [31:0] R10002;
  wire [31:0] R10001;
  wire [31:0] R10000;
  wire [31:0] R9999;
  wire [31:0] R9998;
  wire [31:0] R9997;
  wire [31:0] R9996;
  wire [31:0] R9995;
  wire [31:0] R9994;
  wire [31:0] R9993;
  wire [31:0] R9992;
  wire [31:0] R9991;
  wire [31:0] R9990;
  wire [31:0] R9989;
  wire [31:0] R9988;
  wire [31:0] R9987;
  wire [31:0] R9986;
  wire [31:0] R9985;
  wire [31:0] R9984;
  wire [31:0] R9983;
  wire [31:0] R9982;
  wire [31:0] R9981;
  wire [31:0] R9980;
  wire [31:0] R9979;
  wire [31:0] R9978;
  wire [31:0] R9977;
  wire [31:0] R9976;
  wire [31:0] R9975;
  wire [31:0] R9974;
  wire [63:0] R9973;
  wire [63:0] R9972;
  wire [63:0] R9971;
  wire [31:0] R9970;
  wire [31:0] R9969;
  wire [31:0] R9968;
  wire [31:0] R9967;
  wire [31:0] R9966;
  wire [31:0] R9965;
  wire [31:0] R9964;
  wire [31:0] R9963;
  wire [31:0] R9962;
  wire [31:0] R9961;
  wire [31:0] R9960;
  wire [31:0] R9959;
  wire [31:0] R9958;
  wire [31:0] R9957;
  wire [31:0] R9956;
  wire [31:0] R9955;
  wire [31:0] R9954;
  wire [31:0] R9953;
  wire [31:0] R9952;
  wire [31:0] R9951;
  wire [31:0] R9950;
  wire [31:0] R9949;
  wire [31:0] R9948;
  wire [31:0] R9947;
  wire [31:0] R9946;
  wire [31:0] R9945;
  wire [31:0] R9944;
  wire [31:0] R9943;
  wire [31:0] R9942;
  wire [31:0] R9941;
  wire [31:0] R9940;
  wire [31:0] R9939;
  wire [31:0] R9938;
  wire [31:0] R9937;
  wire [31:0] R9936;
  wire [31:0] R9935;
  wire [31:0] R9934;
  wire [31:0] R9933;
  wire [31:0] R9932;
  wire [31:0] R9931;
  wire [31:0] R9930;
  wire [31:0] R9929;
  wire [31:0] R9928;
  wire [31:0] R9927;
  wire [31:0] R9926;
  wire [31:0] R9925;
  wire [31:0] R9924;
  wire [31:0] R9923;
  wire [31:0] R9922;
  wire [31:0] R9921;
  wire [31:0] R9920;
  wire [31:0] R9919;
  wire [31:0] R9918;
  wire [31:0] R9917;
  wire [31:0] R9916;
  wire [31:0] R9915;
  wire [31:0] R9914;
  wire [31:0] R9913;
  wire [31:0] R9912;
  wire [31:0] R9911;
  wire [31:0] R9910;
  wire [31:0] R9909;
  wire [31:0] R9908;
  wire [31:0] R9907;
  wire [31:0] R9906;
  wire [31:0] R9905;
  wire [31:0] R9904;
  wire [31:0] R9903;
  wire [31:0] R9902;
  wire [31:0] R9901;
  wire [31:0] R9900;
  wire [31:0] R9899;
  wire [31:0] R9898;
  wire [31:0] R9897;
  wire [31:0] R9896;
  wire [31:0] R9895;
  wire [31:0] R9894;
  wire [31:0] R9893;
  wire [31:0] R9892;
  wire [31:0] R9891;
  wire [31:0] R9890;
  wire [31:0] R9889;
  wire [31:0] R9888;
  wire [31:0] R9887;
  wire [31:0] R9886;
  wire [31:0] R9885;
  wire [31:0] R9884;
  wire [31:0] R9883;
  wire [31:0] R9882;
  wire [31:0] R9881;
  wire [31:0] R9880;
  wire [31:0] R9879;
  wire [31:0] R9878;
  wire [31:0] R9877;
  wire [31:0] R9876;
  wire [31:0] R9875;
  wire [31:0] R9874;
  wire [31:0] R9873;
  wire [31:0] R9872;
  wire [31:0] R9871;
  wire [31:0] R9870;
  wire [31:0] R9869;
  wire [31:0] R9868;
  wire [31:0] R9867;
  wire [31:0] R9866;
  wire [31:0] R9865;
  wire [31:0] R9864;
  wire [31:0] R9863;
  wire [31:0] R9862;
  wire [31:0] R9861;
  wire [31:0] R9860;
  wire [31:0] R9859;
  wire [31:0] R9858;
  wire [31:0] R9857;
  wire [31:0] R9856;
  wire [31:0] R9855;
  wire [31:0] R9854;
  wire [31:0] R9853;
  wire [31:0] R9852;
  wire [31:0] R9851;
  wire [31:0] R9850;
  wire [31:0] R9849;
  wire [31:0] R9848;
  wire [31:0] R9847;
  wire [31:0] R9846;
  wire [31:0] R9845;
  wire [31:0] R9844;
  wire [31:0] R9843;
  wire [63:0] R9842;
  wire [31:0] R9841;
  wire [63:0] R9840;
  wire [63:0] R9839;
  wire [63:0] R9838;
  wire [63:0] R9837;
  wire [63:0] R9836;
  wire [63:0] R9835;
  wire [63:0] R9834;
  wire [63:0] R9833;
  wire [63:0] R9832;
  wire [63:0] R9831;
  wire [63:0] R9830;
  wire [63:0] R9829;
  wire [63:0] R9828;
  wire [63:0] R9827;
  wire [63:0] R9826;
  wire [63:0] R9825;
  wire [63:0] R9824;
  wire [63:0] R9823;
  wire [63:0] R9822;
  wire [63:0] R9821;
  wire [63:0] R9820;
  wire [63:0] R9819;
  wire [63:0] R9818;
  wire [63:0] R9817;
  wire [63:0] R9816;
  wire [63:0] R9815;
  wire [63:0] R9814;
  wire [63:0] R9813;
  wire [63:0] R9812;
  wire [63:0] R9811;
  wire [63:0] R9810;
  wire [63:0] R9809;
  wire [63:0] R9808;
  wire [63:0] R9807;
  wire [63:0] R9806;
  wire [63:0] R9805;
  wire [63:0] R9804;
  wire [63:0] R9803;
  wire [63:0] R9802;
  wire [63:0] R9801;
  wire [63:0] R9800;
  wire [63:0] R9799;
  wire [63:0] R9798;
  wire [63:0] R9797;
  wire [63:0] R9796;
  wire [63:0] R9795;
  wire [0:0] R9794;
  wire [0:0] R9793;
  wire [0:0] R9792;
  wire [0:0] R9791;
  wire [0:0] R9790;
  wire [0:0] R9789;
  wire [0:0] R9788;
  wire [0:0] R9787;
  wire [0:0] R9786;
  wire [0:0] R9785;
  wire [0:0] R9784;
  wire [0:0] R9783;
  wire [0:0] R9782;
  wire [0:0] R9781;
  wire [0:0] R9780;
  wire [0:0] R9779;
  wire [0:0] R9778;
  wire [0:0] R9777;
  wire [0:0] R9776;
  wire [0:0] R9775;
  wire [0:0] R9774;
  wire [0:0] R9773;
  wire [0:0] R9772;
  wire [0:0] R9771;
  wire [0:0] R9770;
  wire [0:0] R9769;
  wire [0:0] R9768;
  wire [0:0] R9767;
  wire [0:0] R9766;
  wire [0:0] R9765;
  wire [0:0] R9764;
  wire [0:0] R9763;
  wire [0:0] R9762;
  wire [0:0] R9761;
  wire [0:0] R9760;
  wire [0:0] R9759;
  wire [0:0] R9758;
  wire [0:0] R9757;
  wire [0:0] R9756;
  wire [0:0] R9755;
  wire [0:0] R9754;
  wire [0:0] R9753;
  wire [0:0] R9752;
  wire [0:0] R9751;
  wire [0:0] R9750;
  wire [0:0] R9749;
  wire [0:0] R9748;
  wire [0:0] R9747;
  wire [0:0] R9746;
  wire [0:0] R9745;
  wire [0:0] R9744;
  wire [0:0] R9743;
  wire [0:0] R9742;
  wire [0:0] R9741;
  wire [0:0] R9740;
  wire [0:0] R9739;
  wire [0:0] R9738;
  wire [0:0] R9737;
  wire [0:0] R9736;
  wire [0:0] R9735;
  wire [0:0] R9734;
  wire [0:0] R9733;
  wire [0:0] R9732;
  wire [0:0] R9731;
  wire [0:0] R9730;
  wire [0:0] R9729;
  wire [0:0] R9728;
  wire [0:0] R9727;
  wire [0:0] R9726;
  wire [0:0] R9725;
  wire [0:0] R9724;
  wire [0:0] R9723;
  wire [0:0] R9722;
  wire [0:0] R9721;
  wire [0:0] R9720;
  wire [0:0] R9719;
  wire [0:0] R9718;
  wire [0:0] R9717;
  wire [0:0] R9716;
  wire [0:0] R9715;
  wire [0:0] R9714;
  wire [0:0] R9713;
  wire [0:0] R9712;
  wire [0:0] R9711;
  wire [0:0] R9710;
  wire [0:0] R9709;
  wire [0:0] R9708;
  wire [0:0] R9707;
  wire [0:0] R9706;
  wire [0:0] R9705;
  wire [0:0] R9704;
  wire [0:0] R9703;
  wire [0:0] R9702;
  wire [0:0] R9701;
  wire [0:0] R9700;
  wire [0:0] R9699;
  wire [0:0] R9698;
  wire [0:0] R9697;
  wire [0:0] R9696;
  wire [0:0] R9695;
  wire [0:0] R9694;
  wire [0:0] R9693;
  wire [0:0] R9692;
  wire [0:0] R9691;
  wire [0:0] R9690;
  wire [0:0] R9689;
  wire [0:0] R9688;
  wire [0:0] R9687;
  wire [0:0] R9686;
  wire [0:0] R9685;
  wire [0:0] R9684;
  wire [0:0] R9683;
  wire [0:0] R9682;
  wire [0:0] R9681;
  wire [0:0] R9680;
  wire [0:0] R9679;
  wire [0:0] R9678;
  wire [0:0] R9677;
  wire [0:0] R9676;
  wire [0:0] R9675;
  wire [0:0] R9674;
  wire [0:0] R9673;
  wire [0:0] R9672;
  wire [0:0] R9671;
  wire [0:0] R9670;
  wire [0:0] R9669;
  wire [0:0] R9668;
  wire [0:0] R9667;
  wire [0:0] R9666;
  wire [0:0] R9665;
  wire [0:0] R9664;
  wire [0:0] R9663;
  wire [0:0] R9662;
  wire [0:0] R9661;
  wire [0:0] R9660;
  wire [0:0] R9659;
  wire [0:0] R9658;
  wire [0:0] R9657;
  wire [0:0] R9656;
  wire [0:0] R9655;
  wire [0:0] R9654;
  wire [0:0] R9653;
  wire [63:0] R9652;
  wire [31:0] R9651;
  wire [31:0] R9650;
  wire [31:0] R9649;
  wire [31:0] R9648;
  wire [31:0] R9647;
  wire [31:0] R9646;
  wire [31:0] R9645;
  wire [31:0] R9644;
  wire [31:0] R9643;
  wire [31:0] R9642;
  wire [31:0] R9641;
  wire [31:0] R9640;
  wire [31:0] R9639;
  wire [31:0] R9638;
  wire [31:0] R9637;
  wire [31:0] R9636;
  wire [31:0] R9635;
  wire [31:0] R9634;
  wire [31:0] R9633;
  wire [31:0] R9632;
  wire [31:0] R9631;
  wire [31:0] R9630;
  wire [31:0] R9629;
  wire [31:0] R9628;
  wire [31:0] R9627;
  wire [31:0] R9626;
  wire [31:0] R9625;
  wire [31:0] R9624;
  wire [31:0] R9623;
  wire [31:0] R9622;
  wire [31:0] R9621;
  wire [31:0] R9620;
  wire [31:0] R9619;
  wire [31:0] R9618;
  wire [31:0] R9617;
  wire [31:0] R9616;
  wire [31:0] R9615;
  wire [31:0] R9614;
  wire [31:0] R9613;
  wire [31:0] R9612;
  wire [31:0] R9611;
  wire [31:0] R9610;
  wire [31:0] R9609;
  wire [31:0] R9608;
  wire [31:0] R9607;
  wire [31:0] R9606;
  wire [31:0] R9605;
  wire [31:0] R9604;
  wire [31:0] R9603;
  wire [31:0] R9602;
  wire [31:0] R9601;
  wire [31:0] R9600;
  wire [31:0] R9599;
  wire [31:0] R9598;
  wire [31:0] R9597;
  wire [31:0] R9596;
  wire [31:0] R9595;
  wire [31:0] R9594;
  wire [31:0] R9593;
  wire [31:0] R9592;
  wire [31:0] R9591;
  wire [31:0] R9590;
  wire [31:0] R9589;
  wire [31:0] R9588;
  wire [31:0] R9587;
  wire [31:0] R9586;
  wire [31:0] R9585;
  wire [31:0] R9584;
  wire [31:0] R9583;
  wire [31:0] R9582;
  wire [31:0] R9581;
  wire [31:0] R9580;
  wire [31:0] R9579;
  wire [31:0] R9578;
  wire [31:0] R9577;
  wire [31:0] R9576;
  wire [31:0] R9575;
  wire [31:0] R9574;
  wire [31:0] R9573;
  wire [31:0] R9572;
  wire [31:0] R9571;
  wire [31:0] R9570;
  wire [31:0] R9569;
  wire [31:0] R9568;
  wire [31:0] R9567;
  wire [31:0] R9566;
  wire [31:0] R9565;
  wire [31:0] R9564;
  wire [31:0] R9563;
  wire [31:0] R9562;
  wire [31:0] R9561;
  wire [31:0] R9560;
  wire [31:0] R9559;
  wire [31:0] R9558;
  wire [31:0] R9557;
  wire [31:0] R9556;
  wire [31:0] R9555;
  wire [31:0] R9554;
  wire [31:0] R9553;
  wire [31:0] R9552;
  wire [31:0] R9551;
  wire [31:0] R9550;
  wire [31:0] R9549;
  wire [31:0] R9548;
  wire [31:0] R9547;
  wire [31:0] R9546;
  wire [31:0] R9545;
  wire [31:0] R9544;
  wire [31:0] R9543;
  wire [31:0] R9542;
  wire [31:0] R9541;
  wire [31:0] R9540;
  wire [31:0] R9539;
  wire [31:0] R9538;
  wire [31:0] R9537;
  wire [31:0] R9536;
  wire [31:0] R9535;
  wire [31:0] R9534;
  wire [31:0] R9533;
  wire [31:0] R9532;
  wire [31:0] R9531;
  wire [31:0] R9530;
  wire [31:0] R9529;
  wire [31:0] R9528;
  wire [31:0] R9527;
  wire [31:0] R9526;
  wire [31:0] R9525;
  wire [31:0] R9524;
  wire [31:0] R9523;
  wire [31:0] R9522;
  wire [31:0] R9521;
  wire [31:0] R9520;
  wire [31:0] R9519;
  wire [31:0] R9518;
  wire [31:0] R9517;
  wire [63:0] R9516;
  wire [63:0] R9515;
  wire [63:0] R9514;
  wire [31:0] R9513;
  wire [31:0] R9512;
  wire [31:0] R9511;
  wire [31:0] R9510;
  wire [31:0] R9509;
  wire [31:0] R9508;
  wire [31:0] R9507;
  wire [31:0] R9506;
  wire [31:0] R9505;
  wire [31:0] R9504;
  wire [31:0] R9503;
  wire [31:0] R9502;
  wire [31:0] R9501;
  wire [31:0] R9500;
  wire [31:0] R9499;
  wire [31:0] R9498;
  wire [31:0] R9497;
  wire [31:0] R9496;
  wire [31:0] R9495;
  wire [31:0] R9494;
  wire [31:0] R9493;
  wire [31:0] R9492;
  wire [31:0] R9491;
  wire [31:0] R9490;
  wire [31:0] R9489;
  wire [31:0] R9488;
  wire [31:0] R9487;
  wire [31:0] R9486;
  wire [31:0] R9485;
  wire [31:0] R9484;
  wire [31:0] R9483;
  wire [31:0] R9482;
  wire [31:0] R9481;
  wire [31:0] R9480;
  wire [31:0] R9479;
  wire [31:0] R9478;
  wire [31:0] R9477;
  wire [31:0] R9476;
  wire [31:0] R9475;
  wire [31:0] R9474;
  wire [31:0] R9473;
  wire [31:0] R9472;
  wire [31:0] R9471;
  wire [31:0] R9470;
  wire [31:0] R9469;
  wire [31:0] R9468;
  wire [31:0] R9467;
  wire [31:0] R9466;
  wire [31:0] R9465;
  wire [31:0] R9464;
  wire [31:0] R9463;
  wire [31:0] R9462;
  wire [31:0] R9461;
  wire [31:0] R9460;
  wire [31:0] R9459;
  wire [31:0] R9458;
  wire [31:0] R9457;
  wire [31:0] R9456;
  wire [31:0] R9455;
  wire [31:0] R9454;
  wire [31:0] R9453;
  wire [31:0] R9452;
  wire [31:0] R9451;
  wire [31:0] R9450;
  wire [31:0] R9449;
  wire [31:0] R9448;
  wire [31:0] R9447;
  wire [31:0] R9446;
  wire [31:0] R9445;
  wire [31:0] R9444;
  wire [31:0] R9443;
  wire [31:0] R9442;
  wire [31:0] R9441;
  wire [31:0] R9440;
  wire [31:0] R9439;
  wire [31:0] R9438;
  wire [31:0] R9437;
  wire [31:0] R9436;
  wire [31:0] R9435;
  wire [31:0] R9434;
  wire [31:0] R9433;
  wire [31:0] R9432;
  wire [31:0] R9431;
  wire [31:0] R9430;
  wire [31:0] R9429;
  wire [31:0] R9428;
  wire [31:0] R9427;
  wire [31:0] R9426;
  wire [31:0] R9425;
  wire [31:0] R9424;
  wire [31:0] R9423;
  wire [31:0] R9422;
  wire [31:0] R9421;
  wire [31:0] R9420;
  wire [31:0] R9419;
  wire [31:0] R9418;
  wire [31:0] R9417;
  wire [31:0] R9416;
  wire [31:0] R9415;
  wire [31:0] R9414;
  wire [31:0] R9413;
  wire [31:0] R9412;
  wire [31:0] R9411;
  wire [31:0] R9410;
  wire [31:0] R9409;
  wire [31:0] R9408;
  wire [31:0] R9407;
  wire [31:0] R9406;
  wire [31:0] R9405;
  wire [31:0] R9404;
  wire [31:0] R9403;
  wire [31:0] R9402;
  wire [31:0] R9401;
  wire [31:0] R9400;
  wire [31:0] R9399;
  wire [31:0] R9398;
  wire [31:0] R9397;
  wire [31:0] R9396;
  wire [31:0] R9395;
  wire [31:0] R9394;
  wire [31:0] R9393;
  wire [31:0] R9392;
  wire [31:0] R9391;
  wire [31:0] R9390;
  wire [31:0] R9389;
  wire [31:0] R9388;
  wire [31:0] R9387;
  wire [31:0] R9386;
  wire [31:0] R9385;
  wire [31:0] R9384;
  wire [31:0] R9383;
  wire [31:0] R9382;
  wire [31:0] R9381;
  wire [31:0] R9380;
  wire [31:0] R9379;
  wire [31:0] R9378;
  wire [31:0] R9377;
  wire [31:0] R9376;
  wire [31:0] R9375;
  wire [31:0] R9374;
  wire [31:0] R9373;
  wire [63:0] R9372;
  wire [31:0] R9371;
  wire [63:0] R9370;
  wire [63:0] R9369;
  wire [63:0] R9368;
  wire [63:0] R9367;
  wire [63:0] R9366;
  wire [63:0] R9365;
  wire [63:0] R9364;
  wire [63:0] R9363;
  wire [63:0] R9362;
  wire [63:0] R9361;
  wire [63:0] R9360;
  wire [63:0] R9359;
  wire [63:0] R9358;
  wire [63:0] R9357;
  wire [63:0] R9356;
  wire [63:0] R9355;
  wire [63:0] R9354;
  wire [63:0] R9353;
  wire [63:0] R9352;
  wire [63:0] R9351;
  wire [63:0] R9350;
  wire [63:0] R9349;
  wire [63:0] R9348;
  wire [63:0] R9347;
  wire [63:0] R9346;
  wire [63:0] R9345;
  wire [63:0] R9344;
  wire [63:0] R9343;
  wire [63:0] R9342;
  wire [63:0] R9341;
  wire [63:0] R9340;
  wire [63:0] R9339;
  wire [63:0] R9338;
  wire [63:0] R9337;
  wire [63:0] R9336;
  wire [63:0] R9335;
  wire [63:0] R9334;
  wire [63:0] R9333;
  wire [63:0] R9332;
  wire [63:0] R9331;
  wire [63:0] R9330;
  wire [63:0] R9329;
  wire [63:0] R9328;
  wire [63:0] R9327;
  wire [63:0] R9326;
  wire [63:0] R9325;
  wire [0:0] R9324;
  wire [0:0] R9323;
  wire [0:0] R9322;
  wire [0:0] R9321;
  wire [0:0] R9320;
  wire [0:0] R9319;
  wire [0:0] R9318;
  wire [0:0] R9317;
  wire [0:0] R9316;
  wire [0:0] R9315;
  wire [0:0] R9314;
  wire [0:0] R9313;
  wire [0:0] R9312;
  wire [0:0] R9311;
  wire [0:0] R9310;
  wire [0:0] R9309;
  wire [0:0] R9308;
  wire [0:0] R9307;
  wire [0:0] R9306;
  wire [0:0] R9305;
  wire [0:0] R9304;
  wire [0:0] R9303;
  wire [0:0] R9302;
  wire [0:0] R9301;
  wire [0:0] R9300;
  wire [0:0] R9299;
  wire [0:0] R9298;
  wire [0:0] R9297;
  wire [0:0] R9296;
  wire [0:0] R9295;
  wire [0:0] R9294;
  wire [0:0] R9293;
  wire [0:0] R9292;
  wire [0:0] R9291;
  wire [0:0] R9290;
  wire [0:0] R9289;
  wire [0:0] R9288;
  wire [0:0] R9287;
  wire [0:0] R9286;
  wire [0:0] R9285;
  wire [0:0] R9284;
  wire [0:0] R9283;
  wire [0:0] R9282;
  wire [0:0] R9281;
  wire [0:0] R9280;
  wire [0:0] R9279;
  wire [0:0] R9278;
  wire [0:0] R9277;
  wire [0:0] R9276;
  wire [0:0] R9275;
  wire [0:0] R9274;
  wire [0:0] R9273;
  wire [0:0] R9272;
  wire [0:0] R9271;
  wire [0:0] R9270;
  wire [0:0] R9269;
  wire [0:0] R9268;
  wire [0:0] R9267;
  wire [0:0] R9266;
  wire [0:0] R9265;
  wire [0:0] R9264;
  wire [0:0] R9263;
  wire [0:0] R9262;
  wire [0:0] R9261;
  wire [0:0] R9260;
  wire [0:0] R9259;
  wire [0:0] R9258;
  wire [0:0] R9257;
  wire [0:0] R9256;
  wire [0:0] R9255;
  wire [0:0] R9254;
  wire [0:0] R9253;
  wire [0:0] R9252;
  wire [0:0] R9251;
  wire [0:0] R9250;
  wire [0:0] R9249;
  wire [0:0] R9248;
  wire [0:0] R9247;
  wire [0:0] R9246;
  wire [0:0] R9245;
  wire [0:0] R9244;
  wire [0:0] R9243;
  wire [0:0] R9242;
  wire [0:0] R9241;
  wire [0:0] R9240;
  wire [0:0] R9239;
  wire [0:0] R9238;
  wire [0:0] R9237;
  wire [0:0] R9236;
  wire [0:0] R9235;
  wire [0:0] R9234;
  wire [0:0] R9233;
  wire [0:0] R9232;
  wire [0:0] R9231;
  wire [0:0] R9230;
  wire [0:0] R9229;
  wire [0:0] R9228;
  wire [0:0] R9227;
  wire [0:0] R9226;
  wire [0:0] R9225;
  wire [0:0] R9224;
  wire [0:0] R9223;
  wire [0:0] R9222;
  wire [0:0] R9221;
  wire [0:0] R9220;
  wire [0:0] R9219;
  wire [0:0] R9218;
  wire [0:0] R9217;
  wire [0:0] R9216;
  wire [0:0] R9215;
  wire [0:0] R9214;
  wire [0:0] R9213;
  wire [0:0] R9212;
  wire [0:0] R9211;
  wire [0:0] R9210;
  wire [0:0] R9209;
  wire [0:0] R9208;
  wire [0:0] R9207;
  wire [0:0] R9206;
  wire [0:0] R9205;
  wire [0:0] R9204;
  wire [0:0] R9203;
  wire [0:0] R9202;
  wire [0:0] R9201;
  wire [0:0] R9200;
  wire [0:0] R9199;
  wire [0:0] R9198;
  wire [0:0] R9197;
  wire [0:0] R9196;
  wire [0:0] R9195;
  wire [0:0] R9194;
  wire [0:0] R9193;
  wire [0:0] R9192;
  wire [0:0] R9191;
  wire [0:0] R9190;
  wire [0:0] R9189;
  wire [0:0] R9188;
  wire [0:0] R9187;
  wire [0:0] R9186;
  wire [0:0] R9185;
  wire [0:0] R9184;
  wire [0:0] R9183;
  wire [0:0] R9182;
  wire [0:0] R9181;
  wire [0:0] R9180;
  wire [0:0] R9179;
  wire [0:0] R9178;
  wire [0:0] R9177;
  wire [0:0] R9176;
  wire [0:0] R9175;
  wire [0:0] R9174;
  wire [0:0] R9173;
  wire [0:0] R9172;
  wire [0:0] R9171;
  wire [0:0] R9170;
  wire [63:0] R9169;
  wire [31:0] R9168;
  wire [31:0] R9167;
  wire [31:0] R9166;
  wire [31:0] R9165;
  wire [31:0] R9164;
  wire [31:0] R9163;
  wire [31:0] R9162;
  wire [31:0] R9161;
  wire [31:0] R9160;
  wire [31:0] R9159;
  wire [31:0] R9158;
  wire [31:0] R9157;
  wire [31:0] R9156;
  wire [31:0] R9155;
  wire [31:0] R9154;
  wire [31:0] R9153;
  wire [31:0] R9152;
  wire [31:0] R9151;
  wire [31:0] R9150;
  wire [31:0] R9149;
  wire [31:0] R9148;
  wire [31:0] R9147;
  wire [31:0] R9146;
  wire [31:0] R9145;
  wire [31:0] R9144;
  wire [31:0] R9143;
  wire [31:0] R9142;
  wire [31:0] R9141;
  wire [31:0] R9140;
  wire [31:0] R9139;
  wire [31:0] R9138;
  wire [31:0] R9137;
  wire [31:0] R9136;
  wire [31:0] R9135;
  wire [31:0] R9134;
  wire [31:0] R9133;
  wire [31:0] R9132;
  wire [31:0] R9131;
  wire [31:0] R9130;
  wire [31:0] R9129;
  wire [31:0] R9128;
  wire [31:0] R9127;
  wire [31:0] R9126;
  wire [31:0] R9125;
  wire [31:0] R9124;
  wire [31:0] R9123;
  wire [31:0] R9122;
  wire [31:0] R9121;
  wire [31:0] R9120;
  wire [31:0] R9119;
  wire [31:0] R9118;
  wire [31:0] R9117;
  wire [31:0] R9116;
  wire [31:0] R9115;
  wire [31:0] R9114;
  wire [31:0] R9113;
  wire [31:0] R9112;
  wire [31:0] R9111;
  wire [31:0] R9110;
  wire [31:0] R9109;
  wire [31:0] R9108;
  wire [31:0] R9107;
  wire [31:0] R9106;
  wire [31:0] R9105;
  wire [31:0] R9104;
  wire [31:0] R9103;
  wire [31:0] R9102;
  wire [31:0] R9101;
  wire [31:0] R9100;
  wire [31:0] R9099;
  wire [31:0] R9098;
  wire [31:0] R9097;
  wire [31:0] R9096;
  wire [31:0] R9095;
  wire [31:0] R9094;
  wire [31:0] R9093;
  wire [31:0] R9092;
  wire [31:0] R9091;
  wire [31:0] R9090;
  wire [31:0] R9089;
  wire [31:0] R9088;
  wire [31:0] R9087;
  wire [31:0] R9086;
  wire [31:0] R9085;
  wire [31:0] R9084;
  wire [31:0] R9083;
  wire [31:0] R9082;
  wire [31:0] R9081;
  wire [31:0] R9080;
  wire [31:0] R9079;
  wire [31:0] R9078;
  wire [31:0] R9077;
  wire [31:0] R9076;
  wire [31:0] R9075;
  wire [31:0] R9074;
  wire [31:0] R9073;
  wire [31:0] R9072;
  wire [31:0] R9071;
  wire [31:0] R9070;
  wire [31:0] R9069;
  wire [31:0] R9068;
  wire [31:0] R9067;
  wire [31:0] R9066;
  wire [31:0] R9065;
  wire [31:0] R9064;
  wire [31:0] R9063;
  wire [31:0] R9062;
  wire [31:0] R9061;
  wire [31:0] R9060;
  wire [31:0] R9059;
  wire [31:0] R9058;
  wire [31:0] R9057;
  wire [31:0] R9056;
  wire [31:0] R9055;
  wire [31:0] R9054;
  wire [31:0] R9053;
  wire [31:0] R9052;
  wire [31:0] R9051;
  wire [31:0] R9050;
  wire [31:0] R9049;
  wire [31:0] R9048;
  wire [31:0] R9047;
  wire [31:0] R9046;
  wire [31:0] R9045;
  wire [31:0] R9044;
  wire [31:0] R9043;
  wire [31:0] R9042;
  wire [31:0] R9041;
  wire [31:0] R9040;
  wire [31:0] R9039;
  wire [31:0] R9038;
  wire [31:0] R9037;
  wire [31:0] R9036;
  wire [31:0] R9035;
  wire [31:0] R9034;
  wire [31:0] R9033;
  wire [31:0] R9032;
  wire [31:0] R9031;
  wire [31:0] R9030;
  wire [31:0] R9029;
  wire [31:0] R9028;
  wire [31:0] R9027;
  wire [31:0] R9026;
  wire [31:0] R9025;
  wire [31:0] R9024;
  wire [31:0] R9023;
  wire [31:0] R9022;
  wire [31:0] R9021;
  wire [63:0] R9020;
  wire [63:0] R9019;
  wire [63:0] R9018;
  wire [31:0] R9017;
  wire [31:0] R9016;
  wire [31:0] R9015;
  wire [31:0] R9014;
  wire [31:0] R9013;
  wire [31:0] R9012;
  wire [31:0] R9011;
  wire [31:0] R9010;
  wire [31:0] R9009;
  wire [31:0] R9008;
  wire [31:0] R9007;
  wire [31:0] R9006;
  wire [31:0] R9005;
  wire [31:0] R9004;
  wire [31:0] R9003;
  wire [31:0] R9002;
  wire [31:0] R9001;
  wire [31:0] R9000;
  wire [31:0] R8999;
  wire [31:0] R8998;
  wire [31:0] R8997;
  wire [31:0] R8996;
  wire [31:0] R8995;
  wire [31:0] R8994;
  wire [31:0] R8993;
  wire [31:0] R8992;
  wire [31:0] R8991;
  wire [31:0] R8990;
  wire [31:0] R8989;
  wire [31:0] R8988;
  wire [31:0] R8987;
  wire [31:0] R8986;
  wire [31:0] R8985;
  wire [31:0] R8984;
  wire [31:0] R8983;
  wire [31:0] R8982;
  wire [31:0] R8981;
  wire [31:0] R8980;
  wire [31:0] R8979;
  wire [31:0] R8978;
  wire [31:0] R8977;
  wire [31:0] R8976;
  wire [31:0] R8975;
  wire [31:0] R8974;
  wire [31:0] R8973;
  wire [31:0] R8972;
  wire [31:0] R8971;
  wire [31:0] R8970;
  wire [31:0] R8969;
  wire [31:0] R8968;
  wire [31:0] R8967;
  wire [31:0] R8966;
  wire [31:0] R8965;
  wire [31:0] R8964;
  wire [31:0] R8963;
  wire [31:0] R8962;
  wire [31:0] R8961;
  wire [31:0] R8960;
  wire [31:0] R8959;
  wire [31:0] R8958;
  wire [31:0] R8957;
  wire [31:0] R8956;
  wire [31:0] R8955;
  wire [31:0] R8954;
  wire [31:0] R8953;
  wire [31:0] R8952;
  wire [31:0] R8951;
  wire [31:0] R8950;
  wire [31:0] R8949;
  wire [31:0] R8948;
  wire [31:0] R8947;
  wire [31:0] R8946;
  wire [31:0] R8945;
  wire [31:0] R8944;
  wire [31:0] R8943;
  wire [31:0] R8942;
  wire [31:0] R8941;
  wire [31:0] R8940;
  wire [31:0] R8939;
  wire [31:0] R8938;
  wire [31:0] R8937;
  wire [31:0] R8936;
  wire [31:0] R8935;
  wire [31:0] R8934;
  wire [31:0] R8933;
  wire [31:0] R8932;
  wire [31:0] R8931;
  wire [31:0] R8930;
  wire [31:0] R8929;
  wire [31:0] R8928;
  wire [31:0] R8927;
  wire [31:0] R8926;
  wire [31:0] R8925;
  wire [31:0] R8924;
  wire [31:0] R8923;
  wire [31:0] R8922;
  wire [31:0] R8921;
  wire [31:0] R8920;
  wire [31:0] R8919;
  wire [31:0] R8918;
  wire [31:0] R8917;
  wire [31:0] R8916;
  wire [31:0] R8915;
  wire [31:0] R8914;
  wire [31:0] R8913;
  wire [31:0] R8912;
  wire [31:0] R8911;
  wire [31:0] R8910;
  wire [31:0] R8909;
  wire [31:0] R8908;
  wire [31:0] R8907;
  wire [31:0] R8906;
  wire [31:0] R8905;
  wire [31:0] R8904;
  wire [31:0] R8903;
  wire [31:0] R8902;
  wire [31:0] R8901;
  wire [31:0] R8900;
  wire [31:0] R8899;
  wire [31:0] R8898;
  wire [31:0] R8897;
  wire [31:0] R8896;
  wire [31:0] R8895;
  wire [31:0] R8894;
  wire [31:0] R8893;
  wire [31:0] R8892;
  wire [31:0] R8891;
  wire [31:0] R8890;
  wire [31:0] R8889;
  wire [31:0] R8888;
  wire [31:0] R8887;
  wire [31:0] R8886;
  wire [31:0] R8885;
  wire [31:0] R8884;
  wire [31:0] R8883;
  wire [31:0] R8882;
  wire [31:0] R8881;
  wire [31:0] R8880;
  wire [31:0] R8879;
  wire [31:0] R8878;
  wire [31:0] R8877;
  wire [31:0] R8876;
  wire [31:0] R8875;
  wire [31:0] R8874;
  wire [31:0] R8873;
  wire [31:0] R8872;
  wire [31:0] R8871;
  wire [31:0] R8870;
  wire [31:0] R8869;
  wire [31:0] R8868;
  wire [31:0] R8867;
  wire [31:0] R8866;
  wire [31:0] R8865;
  wire [31:0] R8864;
  wire [63:0] R8863;
  wire [31:0] R8862;
  wire [63:0] R8861;
  wire [63:0] R8860;
  wire [63:0] R8859;
  wire [63:0] R8858;
  wire [63:0] R8857;
  wire [63:0] R8856;
  wire [63:0] R8855;
  wire [63:0] R8854;
  wire [63:0] R8853;
  wire [63:0] R8852;
  wire [63:0] R8851;
  wire [63:0] R8850;
  wire [63:0] R8849;
  wire [63:0] R8848;
  wire [63:0] R8847;
  wire [63:0] R8846;
  wire [63:0] R8845;
  wire [63:0] R8844;
  wire [63:0] R8843;
  wire [63:0] R8842;
  wire [63:0] R8841;
  wire [63:0] R8840;
  wire [63:0] R8839;
  wire [63:0] R8838;
  wire [63:0] R8837;
  wire [63:0] R8836;
  wire [63:0] R8835;
  wire [63:0] R8834;
  wire [63:0] R8833;
  wire [63:0] R8832;
  wire [63:0] R8831;
  wire [63:0] R8830;
  wire [63:0] R8829;
  wire [63:0] R8828;
  wire [63:0] R8827;
  wire [63:0] R8826;
  wire [63:0] R8825;
  wire [63:0] R8824;
  wire [63:0] R8823;
  wire [63:0] R8822;
  wire [63:0] R8821;
  wire [63:0] R8820;
  wire [63:0] R8819;
  wire [63:0] R8818;
  wire [63:0] R8817;
  wire [63:0] R8816;
  wire [0:0] R8815;
  wire [0:0] R8814;
  wire [0:0] R8813;
  wire [0:0] R8812;
  wire [0:0] R8811;
  wire [0:0] R8810;
  wire [0:0] R8809;
  wire [0:0] R8808;
  wire [0:0] R8807;
  wire [0:0] R8806;
  wire [0:0] R8805;
  wire [0:0] R8804;
  wire [0:0] R8803;
  wire [0:0] R8802;
  wire [0:0] R8801;
  wire [0:0] R8800;
  wire [0:0] R8799;
  wire [0:0] R8798;
  wire [0:0] R8797;
  wire [0:0] R8796;
  wire [0:0] R8795;
  wire [0:0] R8794;
  wire [0:0] R8793;
  wire [0:0] R8792;
  wire [0:0] R8791;
  wire [0:0] R8790;
  wire [0:0] R8789;
  wire [0:0] R8788;
  wire [0:0] R8787;
  wire [0:0] R8786;
  wire [0:0] R8785;
  wire [0:0] R8784;
  wire [0:0] R8783;
  wire [0:0] R8782;
  wire [0:0] R8781;
  wire [0:0] R8780;
  wire [0:0] R8779;
  wire [0:0] R8778;
  wire [0:0] R8777;
  wire [0:0] R8776;
  wire [0:0] R8775;
  wire [0:0] R8774;
  wire [0:0] R8773;
  wire [0:0] R8772;
  wire [0:0] R8771;
  wire [0:0] R8770;
  wire [0:0] R8769;
  wire [0:0] R8768;
  wire [0:0] R8767;
  wire [0:0] R8766;
  wire [0:0] R8765;
  wire [0:0] R8764;
  wire [0:0] R8763;
  wire [0:0] R8762;
  wire [0:0] R8761;
  wire [0:0] R8760;
  wire [0:0] R8759;
  wire [0:0] R8758;
  wire [0:0] R8757;
  wire [0:0] R8756;
  wire [0:0] R8755;
  wire [0:0] R8754;
  wire [0:0] R8753;
  wire [0:0] R8752;
  wire [0:0] R8751;
  wire [0:0] R8750;
  wire [0:0] R8749;
  wire [0:0] R8748;
  wire [0:0] R8747;
  wire [0:0] R8746;
  wire [0:0] R8745;
  wire [0:0] R8744;
  wire [0:0] R8743;
  wire [0:0] R8742;
  wire [0:0] R8741;
  wire [0:0] R8740;
  wire [0:0] R8739;
  wire [0:0] R8738;
  wire [0:0] R8737;
  wire [0:0] R8736;
  wire [0:0] R8735;
  wire [0:0] R8734;
  wire [0:0] R8733;
  wire [0:0] R8732;
  wire [0:0] R8731;
  wire [0:0] R8730;
  wire [0:0] R8729;
  wire [0:0] R8728;
  wire [0:0] R8727;
  wire [0:0] R8726;
  wire [0:0] R8725;
  wire [0:0] R8724;
  wire [0:0] R8723;
  wire [0:0] R8722;
  wire [0:0] R8721;
  wire [0:0] R8720;
  wire [0:0] R8719;
  wire [0:0] R8718;
  wire [0:0] R8717;
  wire [0:0] R8716;
  wire [0:0] R8715;
  wire [0:0] R8714;
  wire [0:0] R8713;
  wire [0:0] R8712;
  wire [0:0] R8711;
  wire [0:0] R8710;
  wire [0:0] R8709;
  wire [0:0] R8708;
  wire [0:0] R8707;
  wire [0:0] R8706;
  wire [0:0] R8705;
  wire [0:0] R8704;
  wire [0:0] R8703;
  wire [0:0] R8702;
  wire [0:0] R8701;
  wire [0:0] R8700;
  wire [0:0] R8699;
  wire [0:0] R8698;
  wire [0:0] R8697;
  wire [0:0] R8696;
  wire [0:0] R8695;
  wire [0:0] R8694;
  wire [0:0] R8693;
  wire [0:0] R8692;
  wire [0:0] R8691;
  wire [0:0] R8690;
  wire [0:0] R8689;
  wire [0:0] R8688;
  wire [0:0] R8687;
  wire [0:0] R8686;
  wire [0:0] R8685;
  wire [0:0] R8684;
  wire [0:0] R8683;
  wire [0:0] R8682;
  wire [0:0] R8681;
  wire [0:0] R8680;
  wire [0:0] R8679;
  wire [0:0] R8678;
  wire [0:0] R8677;
  wire [0:0] R8676;
  wire [0:0] R8675;
  wire [0:0] R8674;
  wire [0:0] R8673;
  wire [0:0] R8672;
  wire [0:0] R8671;
  wire [0:0] R8670;
  wire [0:0] R8669;
  wire [0:0] R8668;
  wire [0:0] R8667;
  wire [0:0] R8666;
  wire [0:0] R8665;
  wire [0:0] R8664;
  wire [0:0] R8663;
  wire [0:0] R8662;
  wire [0:0] R8661;
  wire [0:0] R8660;
  wire [0:0] R8659;
  wire [0:0] R8658;
  wire [0:0] R8657;
  wire [0:0] R8656;
  wire [0:0] R8655;
  wire [0:0] R8654;
  wire [0:0] R8653;
  wire [0:0] R8652;
  wire [0:0] R8651;
  wire [0:0] R8650;
  wire [0:0] R8649;
  wire [0:0] R8648;
  wire [63:0] R8647;
  wire [31:0] R8646;
  wire [31:0] R8645;
  wire [31:0] R8644;
  wire [31:0] R8643;
  wire [31:0] R8642;
  wire [31:0] R8641;
  wire [31:0] R8640;
  wire [31:0] R8639;
  wire [31:0] R8638;
  wire [31:0] R8637;
  wire [31:0] R8636;
  wire [31:0] R8635;
  wire [31:0] R8634;
  wire [31:0] R8633;
  wire [31:0] R8632;
  wire [31:0] R8631;
  wire [31:0] R8630;
  wire [31:0] R8629;
  wire [31:0] R8628;
  wire [31:0] R8627;
  wire [31:0] R8626;
  wire [31:0] R8625;
  wire [31:0] R8624;
  wire [31:0] R8623;
  wire [31:0] R8622;
  wire [31:0] R8621;
  wire [31:0] R8620;
  wire [31:0] R8619;
  wire [31:0] R8618;
  wire [31:0] R8617;
  wire [31:0] R8616;
  wire [31:0] R8615;
  wire [31:0] R8614;
  wire [31:0] R8613;
  wire [31:0] R8612;
  wire [31:0] R8611;
  wire [31:0] R8610;
  wire [31:0] R8609;
  wire [31:0] R8608;
  wire [31:0] R8607;
  wire [31:0] R8606;
  wire [31:0] R8605;
  wire [31:0] R8604;
  wire [31:0] R8603;
  wire [31:0] R8602;
  wire [31:0] R8601;
  wire [31:0] R8600;
  wire [31:0] R8599;
  wire [31:0] R8598;
  wire [31:0] R8597;
  wire [31:0] R8596;
  wire [31:0] R8595;
  wire [31:0] R8594;
  wire [31:0] R8593;
  wire [31:0] R8592;
  wire [31:0] R8591;
  wire [31:0] R8590;
  wire [31:0] R8589;
  wire [31:0] R8588;
  wire [31:0] R8587;
  wire [31:0] R8586;
  wire [31:0] R8585;
  wire [31:0] R8584;
  wire [31:0] R8583;
  wire [31:0] R8582;
  wire [31:0] R8581;
  wire [31:0] R8580;
  wire [31:0] R8579;
  wire [31:0] R8578;
  wire [31:0] R8577;
  wire [31:0] R8576;
  wire [31:0] R8575;
  wire [31:0] R8574;
  wire [31:0] R8573;
  wire [31:0] R8572;
  wire [31:0] R8571;
  wire [31:0] R8570;
  wire [31:0] R8569;
  wire [31:0] R8568;
  wire [31:0] R8567;
  wire [31:0] R8566;
  wire [31:0] R8565;
  wire [31:0] R8564;
  wire [31:0] R8563;
  wire [31:0] R8562;
  wire [31:0] R8561;
  wire [31:0] R8560;
  wire [31:0] R8559;
  wire [31:0] R8558;
  wire [31:0] R8557;
  wire [31:0] R8556;
  wire [31:0] R8555;
  wire [31:0] R8554;
  wire [31:0] R8553;
  wire [31:0] R8552;
  wire [31:0] R8551;
  wire [31:0] R8550;
  wire [31:0] R8549;
  wire [31:0] R8548;
  wire [31:0] R8547;
  wire [31:0] R8546;
  wire [31:0] R8545;
  wire [31:0] R8544;
  wire [31:0] R8543;
  wire [31:0] R8542;
  wire [31:0] R8541;
  wire [31:0] R8540;
  wire [31:0] R8539;
  wire [31:0] R8538;
  wire [31:0] R8537;
  wire [31:0] R8536;
  wire [31:0] R8535;
  wire [31:0] R8534;
  wire [31:0] R8533;
  wire [31:0] R8532;
  wire [31:0] R8531;
  wire [31:0] R8530;
  wire [31:0] R8529;
  wire [31:0] R8528;
  wire [31:0] R8527;
  wire [31:0] R8526;
  wire [31:0] R8525;
  wire [31:0] R8524;
  wire [31:0] R8523;
  wire [31:0] R8522;
  wire [31:0] R8521;
  wire [31:0] R8520;
  wire [31:0] R8519;
  wire [31:0] R8518;
  wire [31:0] R8517;
  wire [31:0] R8516;
  wire [31:0] R8515;
  wire [31:0] R8514;
  wire [31:0] R8513;
  wire [31:0] R8512;
  wire [31:0] R8511;
  wire [31:0] R8510;
  wire [31:0] R8509;
  wire [31:0] R8508;
  wire [31:0] R8507;
  wire [31:0] R8506;
  wire [31:0] R8505;
  wire [31:0] R8504;
  wire [31:0] R8503;
  wire [31:0] R8502;
  wire [31:0] R8501;
  wire [31:0] R8500;
  wire [31:0] R8499;
  wire [31:0] R8498;
  wire [31:0] R8497;
  wire [31:0] R8496;
  wire [31:0] R8495;
  wire [31:0] R8494;
  wire [31:0] R8493;
  wire [31:0] R8492;
  wire [31:0] R8491;
  wire [31:0] R8490;
  wire [31:0] R8489;
  wire [31:0] R8488;
  wire [31:0] R8487;
  wire [31:0] R8486;
  wire [63:0] R8485;
  wire [63:0] R8484;
  wire [63:0] R8483;
  wire [31:0] R8482;
  wire [31:0] R8481;
  wire [31:0] R8480;
  wire [31:0] R8479;
  wire [31:0] R8478;
  wire [31:0] R8477;
  wire [31:0] R8476;
  wire [31:0] R8475;
  wire [31:0] R8474;
  wire [31:0] R8473;
  wire [31:0] R8472;
  wire [31:0] R8471;
  wire [31:0] R8470;
  wire [31:0] R8469;
  wire [31:0] R8468;
  wire [31:0] R8467;
  wire [31:0] R8466;
  wire [31:0] R8465;
  wire [31:0] R8464;
  wire [31:0] R8463;
  wire [31:0] R8462;
  wire [31:0] R8461;
  wire [31:0] R8460;
  wire [31:0] R8459;
  wire [31:0] R8458;
  wire [31:0] R8457;
  wire [31:0] R8456;
  wire [31:0] R8455;
  wire [31:0] R8454;
  wire [31:0] R8453;
  wire [31:0] R8452;
  wire [31:0] R8451;
  wire [31:0] R8450;
  wire [31:0] R8449;
  wire [31:0] R8448;
  wire [31:0] R8447;
  wire [31:0] R8446;
  wire [31:0] R8445;
  wire [31:0] R8444;
  wire [31:0] R8443;
  wire [31:0] R8442;
  wire [31:0] R8441;
  wire [31:0] R8440;
  wire [31:0] R8439;
  wire [31:0] R8438;
  wire [31:0] R8437;
  wire [31:0] R8436;
  wire [31:0] R8435;
  wire [31:0] R8434;
  wire [31:0] R8433;
  wire [31:0] R8432;
  wire [31:0] R8431;
  wire [31:0] R8430;
  wire [31:0] R8429;
  wire [31:0] R8428;
  wire [31:0] R8427;
  wire [31:0] R8426;
  wire [31:0] R8425;
  wire [31:0] R8424;
  wire [31:0] R8423;
  wire [31:0] R8422;
  wire [31:0] R8421;
  wire [31:0] R8420;
  wire [31:0] R8419;
  wire [31:0] R8418;
  wire [31:0] R8417;
  wire [31:0] R8416;
  wire [31:0] R8415;
  wire [31:0] R8414;
  wire [31:0] R8413;
  wire [31:0] R8412;
  wire [31:0] R8411;
  wire [31:0] R8410;
  wire [31:0] R8409;
  wire [31:0] R8408;
  wire [31:0] R8407;
  wire [31:0] R8406;
  wire [31:0] R8405;
  wire [31:0] R8404;
  wire [31:0] R8403;
  wire [31:0] R8402;
  wire [31:0] R8401;
  wire [31:0] R8400;
  wire [31:0] R8399;
  wire [31:0] R8398;
  wire [31:0] R8397;
  wire [31:0] R8396;
  wire [31:0] R8395;
  wire [31:0] R8394;
  wire [31:0] R8393;
  wire [31:0] R8392;
  wire [31:0] R8391;
  wire [31:0] R8390;
  wire [31:0] R8389;
  wire [31:0] R8388;
  wire [31:0] R8387;
  wire [31:0] R8386;
  wire [31:0] R8385;
  wire [31:0] R8384;
  wire [31:0] R8383;
  wire [31:0] R8382;
  wire [31:0] R8381;
  wire [31:0] R8380;
  wire [31:0] R8379;
  wire [31:0] R8378;
  wire [31:0] R8377;
  wire [31:0] R8376;
  wire [31:0] R8375;
  wire [31:0] R8374;
  wire [31:0] R8373;
  wire [31:0] R8372;
  wire [31:0] R8371;
  wire [31:0] R8370;
  wire [31:0] R8369;
  wire [31:0] R8368;
  wire [31:0] R8367;
  wire [31:0] R8366;
  wire [31:0] R8365;
  wire [31:0] R8364;
  wire [31:0] R8363;
  wire [31:0] R8362;
  wire [31:0] R8361;
  wire [31:0] R8360;
  wire [31:0] R8359;
  wire [31:0] R8358;
  wire [31:0] R8357;
  wire [31:0] R8356;
  wire [31:0] R8355;
  wire [31:0] R8354;
  wire [31:0] R8353;
  wire [31:0] R8352;
  wire [31:0] R8351;
  wire [31:0] R8350;
  wire [31:0] R8349;
  wire [31:0] R8348;
  wire [31:0] R8347;
  wire [31:0] R8346;
  wire [31:0] R8345;
  wire [31:0] R8344;
  wire [31:0] R8343;
  wire [31:0] R8342;
  wire [31:0] R8341;
  wire [31:0] R8340;
  wire [31:0] R8339;
  wire [31:0] R8338;
  wire [31:0] R8337;
  wire [31:0] R8336;
  wire [31:0] R8335;
  wire [31:0] R8334;
  wire [31:0] R8333;
  wire [31:0] R8332;
  wire [31:0] R8331;
  wire [31:0] R8330;
  wire [31:0] R8329;
  wire [31:0] R8328;
  wire [31:0] R8327;
  wire [31:0] R8326;
  wire [31:0] R8325;
  wire [31:0] R8324;
  wire [31:0] R8323;
  wire [31:0] R8322;
  wire [31:0] R8321;
  wire [31:0] R8320;
  wire [31:0] R8319;
  wire [31:0] R8318;
  wire [31:0] R8317;
  wire [31:0] R8316;
  wire [63:0] R8315;
  wire [31:0] R8314;
  wire [63:0] R8313;
  wire [63:0] R8312;
  wire [63:0] R8311;
  wire [63:0] R8310;
  wire [63:0] R8309;
  wire [63:0] R8308;
  wire [63:0] R8307;
  wire [63:0] R8306;
  wire [63:0] R8305;
  wire [63:0] R8304;
  wire [63:0] R8303;
  wire [63:0] R8302;
  wire [63:0] R8301;
  wire [63:0] R8300;
  wire [63:0] R8299;
  wire [63:0] R8298;
  wire [63:0] R8297;
  wire [63:0] R8296;
  wire [63:0] R8295;
  wire [63:0] R8294;
  wire [63:0] R8293;
  wire [63:0] R8292;
  wire [63:0] R8291;
  wire [63:0] R8290;
  wire [63:0] R8289;
  wire [63:0] R8288;
  wire [63:0] R8287;
  wire [63:0] R8286;
  wire [63:0] R8285;
  wire [63:0] R8284;
  wire [63:0] R8283;
  wire [63:0] R8282;
  wire [63:0] R8281;
  wire [63:0] R8280;
  wire [63:0] R8279;
  wire [63:0] R8278;
  wire [63:0] R8277;
  wire [63:0] R8276;
  wire [63:0] R8275;
  wire [63:0] R8274;
  wire [63:0] R8273;
  wire [63:0] R8272;
  wire [63:0] R8271;
  wire [63:0] R8270;
  wire [63:0] R8269;
  wire [63:0] R8268;
  wire [0:0] R8267;
  wire [0:0] R8266;
  wire [0:0] R8265;
  wire [0:0] R8264;
  wire [0:0] R8263;
  wire [0:0] R8262;
  wire [0:0] R8261;
  wire [0:0] R8260;
  wire [0:0] R8259;
  wire [0:0] R8258;
  wire [0:0] R8257;
  wire [0:0] R8256;
  wire [0:0] R8255;
  wire [0:0] R8254;
  wire [0:0] R8253;
  wire [0:0] R8252;
  wire [0:0] R8251;
  wire [0:0] R8250;
  wire [0:0] R8249;
  wire [0:0] R8248;
  wire [0:0] R8247;
  wire [0:0] R8246;
  wire [0:0] R8245;
  wire [0:0] R8244;
  wire [0:0] R8243;
  wire [0:0] R8242;
  wire [0:0] R8241;
  wire [0:0] R8240;
  wire [0:0] R8239;
  wire [0:0] R8238;
  wire [0:0] R8237;
  wire [0:0] R8236;
  wire [0:0] R8235;
  wire [0:0] R8234;
  wire [0:0] R8233;
  wire [0:0] R8232;
  wire [0:0] R8231;
  wire [0:0] R8230;
  wire [0:0] R8229;
  wire [0:0] R8228;
  wire [0:0] R8227;
  wire [0:0] R8226;
  wire [0:0] R8225;
  wire [0:0] R8224;
  wire [0:0] R8223;
  wire [0:0] R8222;
  wire [0:0] R8221;
  wire [0:0] R8220;
  wire [0:0] R8219;
  wire [0:0] R8218;
  wire [0:0] R8217;
  wire [0:0] R8216;
  wire [0:0] R8215;
  wire [0:0] R8214;
  wire [0:0] R8213;
  wire [0:0] R8212;
  wire [0:0] R8211;
  wire [0:0] R8210;
  wire [0:0] R8209;
  wire [0:0] R8208;
  wire [0:0] R8207;
  wire [0:0] R8206;
  wire [0:0] R8205;
  wire [0:0] R8204;
  wire [0:0] R8203;
  wire [0:0] R8202;
  wire [0:0] R8201;
  wire [0:0] R8200;
  wire [0:0] R8199;
  wire [0:0] R8198;
  wire [0:0] R8197;
  wire [0:0] R8196;
  wire [0:0] R8195;
  wire [0:0] R8194;
  wire [0:0] R8193;
  wire [0:0] R8192;
  wire [0:0] R8191;
  wire [0:0] R8190;
  wire [0:0] R8189;
  wire [0:0] R8188;
  wire [0:0] R8187;
  wire [0:0] R8186;
  wire [0:0] R8185;
  wire [0:0] R8184;
  wire [0:0] R8183;
  wire [0:0] R8182;
  wire [0:0] R8181;
  wire [0:0] R8180;
  wire [0:0] R8179;
  wire [0:0] R8178;
  wire [0:0] R8177;
  wire [0:0] R8176;
  wire [0:0] R8175;
  wire [0:0] R8174;
  wire [0:0] R8173;
  wire [0:0] R8172;
  wire [0:0] R8171;
  wire [0:0] R8170;
  wire [0:0] R8169;
  wire [0:0] R8168;
  wire [0:0] R8167;
  wire [0:0] R8166;
  wire [0:0] R8165;
  wire [0:0] R8164;
  wire [0:0] R8163;
  wire [0:0] R8162;
  wire [0:0] R8161;
  wire [0:0] R8160;
  wire [0:0] R8159;
  wire [0:0] R8158;
  wire [0:0] R8157;
  wire [0:0] R8156;
  wire [0:0] R8155;
  wire [0:0] R8154;
  wire [0:0] R8153;
  wire [0:0] R8152;
  wire [0:0] R8151;
  wire [0:0] R8150;
  wire [0:0] R8149;
  wire [0:0] R8148;
  wire [0:0] R8147;
  wire [0:0] R8146;
  wire [0:0] R8145;
  wire [0:0] R8144;
  wire [0:0] R8143;
  wire [0:0] R8142;
  wire [0:0] R8141;
  wire [0:0] R8140;
  wire [0:0] R8139;
  wire [0:0] R8138;
  wire [0:0] R8137;
  wire [0:0] R8136;
  wire [0:0] R8135;
  wire [0:0] R8134;
  wire [0:0] R8133;
  wire [0:0] R8132;
  wire [0:0] R8131;
  wire [0:0] R8130;
  wire [0:0] R8129;
  wire [0:0] R8128;
  wire [0:0] R8127;
  wire [0:0] R8126;
  wire [0:0] R8125;
  wire [0:0] R8124;
  wire [0:0] R8123;
  wire [0:0] R8122;
  wire [0:0] R8121;
  wire [0:0] R8120;
  wire [0:0] R8119;
  wire [0:0] R8118;
  wire [0:0] R8117;
  wire [0:0] R8116;
  wire [0:0] R8115;
  wire [0:0] R8114;
  wire [0:0] R8113;
  wire [0:0] R8112;
  wire [0:0] R8111;
  wire [0:0] R8110;
  wire [0:0] R8109;
  wire [0:0] R8108;
  wire [0:0] R8107;
  wire [0:0] R8106;
  wire [0:0] R8105;
  wire [0:0] R8104;
  wire [0:0] R8103;
  wire [0:0] R8102;
  wire [0:0] R8101;
  wire [0:0] R8100;
  wire [0:0] R8099;
  wire [0:0] R8098;
  wire [0:0] R8097;
  wire [0:0] R8096;
  wire [0:0] R8095;
  wire [0:0] R8094;
  wire [0:0] R8093;
  wire [0:0] R8092;
  wire [0:0] R8091;
  wire [0:0] R8090;
  wire [0:0] R8089;
  wire [0:0] R8088;
  wire [0:0] R8087;
  wire [63:0] R8086;
  wire [31:0] R8085;
  wire [31:0] R8084;
  wire [31:0] R8083;
  wire [31:0] R8082;
  wire [31:0] R8081;
  wire [31:0] R8080;
  wire [31:0] R8079;
  wire [31:0] R8078;
  wire [31:0] R8077;
  wire [31:0] R8076;
  wire [31:0] R8075;
  wire [31:0] R8074;
  wire [31:0] R8073;
  wire [31:0] R8072;
  wire [31:0] R8071;
  wire [31:0] R8070;
  wire [31:0] R8069;
  wire [31:0] R8068;
  wire [31:0] R8067;
  wire [31:0] R8066;
  wire [31:0] R8065;
  wire [31:0] R8064;
  wire [31:0] R8063;
  wire [31:0] R8062;
  wire [31:0] R8061;
  wire [31:0] R8060;
  wire [31:0] R8059;
  wire [31:0] R8058;
  wire [31:0] R8057;
  wire [31:0] R8056;
  wire [31:0] R8055;
  wire [31:0] R8054;
  wire [31:0] R8053;
  wire [31:0] R8052;
  wire [31:0] R8051;
  wire [31:0] R8050;
  wire [31:0] R8049;
  wire [31:0] R8048;
  wire [31:0] R8047;
  wire [31:0] R8046;
  wire [31:0] R8045;
  wire [31:0] R8044;
  wire [31:0] R8043;
  wire [31:0] R8042;
  wire [31:0] R8041;
  wire [31:0] R8040;
  wire [31:0] R8039;
  wire [31:0] R8038;
  wire [31:0] R8037;
  wire [31:0] R8036;
  wire [31:0] R8035;
  wire [31:0] R8034;
  wire [31:0] R8033;
  wire [31:0] R8032;
  wire [31:0] R8031;
  wire [31:0] R8030;
  wire [31:0] R8029;
  wire [31:0] R8028;
  wire [31:0] R8027;
  wire [31:0] R8026;
  wire [31:0] R8025;
  wire [31:0] R8024;
  wire [31:0] R8023;
  wire [31:0] R8022;
  wire [31:0] R8021;
  wire [31:0] R8020;
  wire [31:0] R8019;
  wire [31:0] R8018;
  wire [31:0] R8017;
  wire [31:0] R8016;
  wire [31:0] R8015;
  wire [31:0] R8014;
  wire [31:0] R8013;
  wire [31:0] R8012;
  wire [31:0] R8011;
  wire [31:0] R8010;
  wire [31:0] R8009;
  wire [31:0] R8008;
  wire [31:0] R8007;
  wire [31:0] R8006;
  wire [31:0] R8005;
  wire [31:0] R8004;
  wire [31:0] R8003;
  wire [31:0] R8002;
  wire [31:0] R8001;
  wire [31:0] R8000;
  wire [31:0] R7999;
  wire [31:0] R7998;
  wire [31:0] R7997;
  wire [31:0] R7996;
  wire [31:0] R7995;
  wire [31:0] R7994;
  wire [31:0] R7993;
  wire [31:0] R7992;
  wire [31:0] R7991;
  wire [31:0] R7990;
  wire [31:0] R7989;
  wire [31:0] R7988;
  wire [31:0] R7987;
  wire [31:0] R7986;
  wire [31:0] R7985;
  wire [31:0] R7984;
  wire [31:0] R7983;
  wire [31:0] R7982;
  wire [31:0] R7981;
  wire [31:0] R7980;
  wire [31:0] R7979;
  wire [31:0] R7978;
  wire [31:0] R7977;
  wire [31:0] R7976;
  wire [31:0] R7975;
  wire [31:0] R7974;
  wire [31:0] R7973;
  wire [31:0] R7972;
  wire [31:0] R7971;
  wire [31:0] R7970;
  wire [31:0] R7969;
  wire [31:0] R7968;
  wire [31:0] R7967;
  wire [31:0] R7966;
  wire [31:0] R7965;
  wire [31:0] R7964;
  wire [31:0] R7963;
  wire [31:0] R7962;
  wire [31:0] R7961;
  wire [31:0] R7960;
  wire [31:0] R7959;
  wire [31:0] R7958;
  wire [31:0] R7957;
  wire [31:0] R7956;
  wire [31:0] R7955;
  wire [31:0] R7954;
  wire [31:0] R7953;
  wire [31:0] R7952;
  wire [31:0] R7951;
  wire [31:0] R7950;
  wire [31:0] R7949;
  wire [31:0] R7948;
  wire [31:0] R7947;
  wire [31:0] R7946;
  wire [31:0] R7945;
  wire [31:0] R7944;
  wire [31:0] R7943;
  wire [31:0] R7942;
  wire [31:0] R7941;
  wire [31:0] R7940;
  wire [31:0] R7939;
  wire [31:0] R7938;
  wire [31:0] R7937;
  wire [31:0] R7936;
  wire [31:0] R7935;
  wire [31:0] R7934;
  wire [31:0] R7933;
  wire [31:0] R7932;
  wire [31:0] R7931;
  wire [31:0] R7930;
  wire [31:0] R7929;
  wire [31:0] R7928;
  wire [31:0] R7927;
  wire [31:0] R7926;
  wire [31:0] R7925;
  wire [31:0] R7924;
  wire [31:0] R7923;
  wire [31:0] R7922;
  wire [31:0] R7921;
  wire [31:0] R7920;
  wire [31:0] R7919;
  wire [31:0] R7918;
  wire [31:0] R7917;
  wire [31:0] R7916;
  wire [31:0] R7915;
  wire [31:0] R7914;
  wire [31:0] R7913;
  wire [31:0] R7912;
  wire [63:0] R7911;
  wire [63:0] R7910;
  wire [63:0] R7909;
  wire [31:0] R7908;
  wire [31:0] R7907;
  wire [31:0] R7906;
  wire [31:0] R7905;
  wire [31:0] R7904;
  wire [31:0] R7903;
  wire [31:0] R7902;
  wire [31:0] R7901;
  wire [31:0] R7900;
  wire [31:0] R7899;
  wire [31:0] R7898;
  wire [31:0] R7897;
  wire [31:0] R7896;
  wire [31:0] R7895;
  wire [31:0] R7894;
  wire [31:0] R7893;
  wire [31:0] R7892;
  wire [31:0] R7891;
  wire [31:0] R7890;
  wire [31:0] R7889;
  wire [31:0] R7888;
  wire [31:0] R7887;
  wire [31:0] R7886;
  wire [31:0] R7885;
  wire [31:0] R7884;
  wire [31:0] R7883;
  wire [31:0] R7882;
  wire [31:0] R7881;
  wire [31:0] R7880;
  wire [31:0] R7879;
  wire [31:0] R7878;
  wire [31:0] R7877;
  wire [31:0] R7876;
  wire [31:0] R7875;
  wire [31:0] R7874;
  wire [31:0] R7873;
  wire [31:0] R7872;
  wire [31:0] R7871;
  wire [31:0] R7870;
  wire [31:0] R7869;
  wire [31:0] R7868;
  wire [31:0] R7867;
  wire [31:0] R7866;
  wire [31:0] R7865;
  wire [31:0] R7864;
  wire [31:0] R7863;
  wire [31:0] R7862;
  wire [31:0] R7861;
  wire [31:0] R7860;
  wire [31:0] R7859;
  wire [31:0] R7858;
  wire [31:0] R7857;
  wire [31:0] R7856;
  wire [31:0] R7855;
  wire [31:0] R7854;
  wire [31:0] R7853;
  wire [31:0] R7852;
  wire [31:0] R7851;
  wire [31:0] R7850;
  wire [31:0] R7849;
  wire [31:0] R7848;
  wire [31:0] R7847;
  wire [31:0] R7846;
  wire [31:0] R7845;
  wire [31:0] R7844;
  wire [31:0] R7843;
  wire [31:0] R7842;
  wire [31:0] R7841;
  wire [31:0] R7840;
  wire [31:0] R7839;
  wire [31:0] R7838;
  wire [31:0] R7837;
  wire [31:0] R7836;
  wire [31:0] R7835;
  wire [31:0] R7834;
  wire [31:0] R7833;
  wire [31:0] R7832;
  wire [31:0] R7831;
  wire [31:0] R7830;
  wire [31:0] R7829;
  wire [31:0] R7828;
  wire [31:0] R7827;
  wire [31:0] R7826;
  wire [31:0] R7825;
  wire [31:0] R7824;
  wire [31:0] R7823;
  wire [31:0] R7822;
  wire [31:0] R7821;
  wire [31:0] R7820;
  wire [31:0] R7819;
  wire [31:0] R7818;
  wire [31:0] R7817;
  wire [31:0] R7816;
  wire [31:0] R7815;
  wire [31:0] R7814;
  wire [31:0] R7813;
  wire [31:0] R7812;
  wire [31:0] R7811;
  wire [31:0] R7810;
  wire [31:0] R7809;
  wire [31:0] R7808;
  wire [31:0] R7807;
  wire [31:0] R7806;
  wire [31:0] R7805;
  wire [31:0] R7804;
  wire [31:0] R7803;
  wire [31:0] R7802;
  wire [31:0] R7801;
  wire [31:0] R7800;
  wire [31:0] R7799;
  wire [31:0] R7798;
  wire [31:0] R7797;
  wire [31:0] R7796;
  wire [31:0] R7795;
  wire [31:0] R7794;
  wire [31:0] R7793;
  wire [31:0] R7792;
  wire [31:0] R7791;
  wire [31:0] R7790;
  wire [31:0] R7789;
  wire [31:0] R7788;
  wire [31:0] R7787;
  wire [31:0] R7786;
  wire [31:0] R7785;
  wire [31:0] R7784;
  wire [31:0] R7783;
  wire [31:0] R7782;
  wire [31:0] R7781;
  wire [31:0] R7780;
  wire [31:0] R7779;
  wire [31:0] R7778;
  wire [31:0] R7777;
  wire [31:0] R7776;
  wire [31:0] R7775;
  wire [31:0] R7774;
  wire [31:0] R7773;
  wire [31:0] R7772;
  wire [31:0] R7771;
  wire [31:0] R7770;
  wire [31:0] R7769;
  wire [31:0] R7768;
  wire [31:0] R7767;
  wire [31:0] R7766;
  wire [31:0] R7765;
  wire [31:0] R7764;
  wire [31:0] R7763;
  wire [31:0] R7762;
  wire [31:0] R7761;
  wire [31:0] R7760;
  wire [31:0] R7759;
  wire [31:0] R7758;
  wire [31:0] R7757;
  wire [31:0] R7756;
  wire [31:0] R7755;
  wire [31:0] R7754;
  wire [31:0] R7753;
  wire [31:0] R7752;
  wire [31:0] R7751;
  wire [31:0] R7750;
  wire [31:0] R7749;
  wire [31:0] R7748;
  wire [31:0] R7747;
  wire [31:0] R7746;
  wire [31:0] R7745;
  wire [31:0] R7744;
  wire [31:0] R7743;
  wire [31:0] R7742;
  wire [31:0] R7741;
  wire [31:0] R7740;
  wire [31:0] R7739;
  wire [31:0] R7738;
  wire [31:0] R7737;
  wire [31:0] R7736;
  wire [31:0] R7735;
  wire [31:0] R7734;
  wire [31:0] R7733;
  wire [31:0] R7732;
  wire [31:0] R7731;
  wire [31:0] R7730;
  wire [31:0] R7729;
  wire [63:0] R7728;
  wire [31:0] R7727;
  wire [63:0] R7726;
  wire [63:0] R7725;
  wire [63:0] R7724;
  wire [63:0] R7723;
  wire [63:0] R7722;
  wire [63:0] R7721;
  wire [63:0] R7720;
  wire [63:0] R7719;
  wire [63:0] R7718;
  wire [63:0] R7717;
  wire [63:0] R7716;
  wire [63:0] R7715;
  wire [63:0] R7714;
  wire [63:0] R7713;
  wire [63:0] R7712;
  wire [63:0] R7711;
  wire [63:0] R7710;
  wire [63:0] R7709;
  wire [63:0] R7708;
  wire [63:0] R7707;
  wire [63:0] R7706;
  wire [63:0] R7705;
  wire [63:0] R7704;
  wire [63:0] R7703;
  wire [63:0] R7702;
  wire [63:0] R7701;
  wire [63:0] R7700;
  wire [63:0] R7699;
  wire [63:0] R7698;
  wire [63:0] R7697;
  wire [63:0] R7696;
  wire [63:0] R7695;
  wire [63:0] R7694;
  wire [63:0] R7693;
  wire [63:0] R7692;
  wire [63:0] R7691;
  wire [63:0] R7690;
  wire [63:0] R7689;
  wire [63:0] R7688;
  wire [63:0] R7687;
  wire [63:0] R7686;
  wire [63:0] R7685;
  wire [63:0] R7684;
  wire [63:0] R7683;
  wire [63:0] R7682;
  wire [63:0] R7681;
  wire [0:0] R7680;
  wire [0:0] R7679;
  wire [0:0] R7678;
  wire [0:0] R7677;
  wire [0:0] R7676;
  wire [0:0] R7675;
  wire [0:0] R7674;
  wire [0:0] R7673;
  wire [0:0] R7672;
  wire [0:0] R7671;
  wire [0:0] R7670;
  wire [0:0] R7669;
  wire [0:0] R7668;
  wire [0:0] R7667;
  wire [0:0] R7666;
  wire [0:0] R7665;
  wire [0:0] R7664;
  wire [0:0] R7663;
  wire [0:0] R7662;
  wire [0:0] R7661;
  wire [0:0] R7660;
  wire [0:0] R7659;
  wire [0:0] R7658;
  wire [0:0] R7657;
  wire [0:0] R7656;
  wire [0:0] R7655;
  wire [0:0] R7654;
  wire [0:0] R7653;
  wire [0:0] R7652;
  wire [0:0] R7651;
  wire [0:0] R7650;
  wire [0:0] R7649;
  wire [0:0] R7648;
  wire [0:0] R7647;
  wire [0:0] R7646;
  wire [0:0] R7645;
  wire [0:0] R7644;
  wire [0:0] R7643;
  wire [0:0] R7642;
  wire [0:0] R7641;
  wire [0:0] R7640;
  wire [0:0] R7639;
  wire [0:0] R7638;
  wire [0:0] R7637;
  wire [0:0] R7636;
  wire [0:0] R7635;
  wire [0:0] R7634;
  wire [0:0] R7633;
  wire [0:0] R7632;
  wire [0:0] R7631;
  wire [0:0] R7630;
  wire [0:0] R7629;
  wire [0:0] R7628;
  wire [0:0] R7627;
  wire [0:0] R7626;
  wire [0:0] R7625;
  wire [0:0] R7624;
  wire [0:0] R7623;
  wire [0:0] R7622;
  wire [0:0] R7621;
  wire [0:0] R7620;
  wire [0:0] R7619;
  wire [0:0] R7618;
  wire [0:0] R7617;
  wire [0:0] R7616;
  wire [0:0] R7615;
  wire [0:0] R7614;
  wire [0:0] R7613;
  wire [0:0] R7612;
  wire [0:0] R7611;
  wire [0:0] R7610;
  wire [0:0] R7609;
  wire [0:0] R7608;
  wire [0:0] R7607;
  wire [0:0] R7606;
  wire [0:0] R7605;
  wire [0:0] R7604;
  wire [0:0] R7603;
  wire [0:0] R7602;
  wire [0:0] R7601;
  wire [0:0] R7600;
  wire [0:0] R7599;
  wire [0:0] R7598;
  wire [0:0] R7597;
  wire [0:0] R7596;
  wire [0:0] R7595;
  wire [0:0] R7594;
  wire [0:0] R7593;
  wire [0:0] R7592;
  wire [0:0] R7591;
  wire [0:0] R7590;
  wire [0:0] R7589;
  wire [0:0] R7588;
  wire [0:0] R7587;
  wire [0:0] R7586;
  wire [0:0] R7585;
  wire [0:0] R7584;
  wire [0:0] R7583;
  wire [0:0] R7582;
  wire [0:0] R7581;
  wire [0:0] R7580;
  wire [0:0] R7579;
  wire [0:0] R7578;
  wire [0:0] R7577;
  wire [0:0] R7576;
  wire [0:0] R7575;
  wire [0:0] R7574;
  wire [0:0] R7573;
  wire [0:0] R7572;
  wire [0:0] R7571;
  wire [0:0] R7570;
  wire [0:0] R7569;
  wire [0:0] R7568;
  wire [0:0] R7567;
  wire [0:0] R7566;
  wire [0:0] R7565;
  wire [0:0] R7564;
  wire [0:0] R7563;
  wire [0:0] R7562;
  wire [0:0] R7561;
  wire [0:0] R7560;
  wire [0:0] R7559;
  wire [0:0] R7558;
  wire [0:0] R7557;
  wire [0:0] R7556;
  wire [0:0] R7555;
  wire [0:0] R7554;
  wire [0:0] R7553;
  wire [0:0] R7552;
  wire [0:0] R7551;
  wire [0:0] R7550;
  wire [0:0] R7549;
  wire [0:0] R7548;
  wire [0:0] R7547;
  wire [0:0] R7546;
  wire [0:0] R7545;
  wire [0:0] R7544;
  wire [0:0] R7543;
  wire [0:0] R7542;
  wire [0:0] R7541;
  wire [0:0] R7540;
  wire [0:0] R7539;
  wire [0:0] R7538;
  wire [0:0] R7537;
  wire [0:0] R7536;
  wire [0:0] R7535;
  wire [0:0] R7534;
  wire [0:0] R7533;
  wire [0:0] R7532;
  wire [0:0] R7531;
  wire [0:0] R7530;
  wire [0:0] R7529;
  wire [0:0] R7528;
  wire [0:0] R7527;
  wire [0:0] R7526;
  wire [0:0] R7525;
  wire [0:0] R7524;
  wire [0:0] R7523;
  wire [0:0] R7522;
  wire [0:0] R7521;
  wire [0:0] R7520;
  wire [0:0] R7519;
  wire [0:0] R7518;
  wire [0:0] R7517;
  wire [0:0] R7516;
  wire [0:0] R7515;
  wire [0:0] R7514;
  wire [0:0] R7513;
  wire [0:0] R7512;
  wire [0:0] R7511;
  wire [0:0] R7510;
  wire [0:0] R7509;
  wire [0:0] R7508;
  wire [0:0] R7507;
  wire [0:0] R7506;
  wire [0:0] R7505;
  wire [0:0] R7504;
  wire [0:0] R7503;
  wire [0:0] R7502;
  wire [0:0] R7501;
  wire [0:0] R7500;
  wire [0:0] R7499;
  wire [0:0] R7498;
  wire [0:0] R7497;
  wire [0:0] R7496;
  wire [0:0] R7495;
  wire [0:0] R7494;
  wire [0:0] R7493;
  wire [0:0] R7492;
  wire [0:0] R7491;
  wire [0:0] R7490;
  wire [0:0] R7489;
  wire [0:0] R7488;
  wire [0:0] R7487;
  wire [63:0] R7486;
  wire [31:0] R7485;
  wire [31:0] R7484;
  wire [31:0] R7483;
  wire [31:0] R7482;
  wire [31:0] R7481;
  wire [31:0] R7480;
  wire [31:0] R7479;
  wire [31:0] R7478;
  wire [31:0] R7477;
  wire [31:0] R7476;
  wire [31:0] R7475;
  wire [31:0] R7474;
  wire [31:0] R7473;
  wire [31:0] R7472;
  wire [31:0] R7471;
  wire [31:0] R7470;
  wire [31:0] R7469;
  wire [31:0] R7468;
  wire [31:0] R7467;
  wire [31:0] R7466;
  wire [31:0] R7465;
  wire [31:0] R7464;
  wire [31:0] R7463;
  wire [31:0] R7462;
  wire [31:0] R7461;
  wire [31:0] R7460;
  wire [31:0] R7459;
  wire [31:0] R7458;
  wire [31:0] R7457;
  wire [31:0] R7456;
  wire [31:0] R7455;
  wire [31:0] R7454;
  wire [31:0] R7453;
  wire [31:0] R7452;
  wire [31:0] R7451;
  wire [31:0] R7450;
  wire [31:0] R7449;
  wire [31:0] R7448;
  wire [31:0] R7447;
  wire [31:0] R7446;
  wire [31:0] R7445;
  wire [31:0] R7444;
  wire [31:0] R7443;
  wire [31:0] R7442;
  wire [31:0] R7441;
  wire [31:0] R7440;
  wire [31:0] R7439;
  wire [31:0] R7438;
  wire [31:0] R7437;
  wire [31:0] R7436;
  wire [31:0] R7435;
  wire [31:0] R7434;
  wire [31:0] R7433;
  wire [31:0] R7432;
  wire [31:0] R7431;
  wire [31:0] R7430;
  wire [31:0] R7429;
  wire [31:0] R7428;
  wire [31:0] R7427;
  wire [31:0] R7426;
  wire [31:0] R7425;
  wire [31:0] R7424;
  wire [31:0] R7423;
  wire [31:0] R7422;
  wire [31:0] R7421;
  wire [31:0] R7420;
  wire [31:0] R7419;
  wire [31:0] R7418;
  wire [31:0] R7417;
  wire [31:0] R7416;
  wire [31:0] R7415;
  wire [31:0] R7414;
  wire [31:0] R7413;
  wire [31:0] R7412;
  wire [31:0] R7411;
  wire [31:0] R7410;
  wire [31:0] R7409;
  wire [31:0] R7408;
  wire [31:0] R7407;
  wire [31:0] R7406;
  wire [31:0] R7405;
  wire [31:0] R7404;
  wire [31:0] R7403;
  wire [31:0] R7402;
  wire [31:0] R7401;
  wire [31:0] R7400;
  wire [31:0] R7399;
  wire [31:0] R7398;
  wire [31:0] R7397;
  wire [31:0] R7396;
  wire [31:0] R7395;
  wire [31:0] R7394;
  wire [31:0] R7393;
  wire [31:0] R7392;
  wire [31:0] R7391;
  wire [31:0] R7390;
  wire [31:0] R7389;
  wire [31:0] R7388;
  wire [31:0] R7387;
  wire [31:0] R7386;
  wire [31:0] R7385;
  wire [31:0] R7384;
  wire [31:0] R7383;
  wire [31:0] R7382;
  wire [31:0] R7381;
  wire [31:0] R7380;
  wire [31:0] R7379;
  wire [31:0] R7378;
  wire [31:0] R7377;
  wire [31:0] R7376;
  wire [31:0] R7375;
  wire [31:0] R7374;
  wire [31:0] R7373;
  wire [31:0] R7372;
  wire [31:0] R7371;
  wire [31:0] R7370;
  wire [31:0] R7369;
  wire [31:0] R7368;
  wire [31:0] R7367;
  wire [31:0] R7366;
  wire [31:0] R7365;
  wire [31:0] R7364;
  wire [31:0] R7363;
  wire [31:0] R7362;
  wire [31:0] R7361;
  wire [31:0] R7360;
  wire [31:0] R7359;
  wire [31:0] R7358;
  wire [31:0] R7357;
  wire [31:0] R7356;
  wire [31:0] R7355;
  wire [31:0] R7354;
  wire [31:0] R7353;
  wire [31:0] R7352;
  wire [31:0] R7351;
  wire [31:0] R7350;
  wire [31:0] R7349;
  wire [31:0] R7348;
  wire [31:0] R7347;
  wire [31:0] R7346;
  wire [31:0] R7345;
  wire [31:0] R7344;
  wire [31:0] R7343;
  wire [31:0] R7342;
  wire [31:0] R7341;
  wire [31:0] R7340;
  wire [31:0] R7339;
  wire [31:0] R7338;
  wire [31:0] R7337;
  wire [31:0] R7336;
  wire [31:0] R7335;
  wire [31:0] R7334;
  wire [31:0] R7333;
  wire [31:0] R7332;
  wire [31:0] R7331;
  wire [31:0] R7330;
  wire [31:0] R7329;
  wire [31:0] R7328;
  wire [31:0] R7327;
  wire [31:0] R7326;
  wire [31:0] R7325;
  wire [31:0] R7324;
  wire [31:0] R7323;
  wire [31:0] R7322;
  wire [31:0] R7321;
  wire [31:0] R7320;
  wire [31:0] R7319;
  wire [31:0] R7318;
  wire [31:0] R7317;
  wire [31:0] R7316;
  wire [31:0] R7315;
  wire [31:0] R7314;
  wire [31:0] R7313;
  wire [31:0] R7312;
  wire [31:0] R7311;
  wire [31:0] R7310;
  wire [31:0] R7309;
  wire [31:0] R7308;
  wire [31:0] R7307;
  wire [31:0] R7306;
  wire [31:0] R7305;
  wire [31:0] R7304;
  wire [31:0] R7303;
  wire [31:0] R7302;
  wire [31:0] R7301;
  wire [31:0] R7300;
  wire [31:0] R7299;
  wire [63:0] R7298;
  wire [63:0] R7297;
  wire [63:0] R7296;
  wire [31:0] R7295;
  wire [31:0] R7294;
  wire [31:0] R7293;
  wire [31:0] R7292;
  wire [31:0] R7291;
  wire [31:0] R7290;
  wire [31:0] R7289;
  wire [31:0] R7288;
  wire [31:0] R7287;
  wire [31:0] R7286;
  wire [31:0] R7285;
  wire [31:0] R7284;
  wire [31:0] R7283;
  wire [31:0] R7282;
  wire [31:0] R7281;
  wire [31:0] R7280;
  wire [31:0] R7279;
  wire [31:0] R7278;
  wire [31:0] R7277;
  wire [31:0] R7276;
  wire [31:0] R7275;
  wire [31:0] R7274;
  wire [31:0] R7273;
  wire [31:0] R7272;
  wire [31:0] R7271;
  wire [31:0] R7270;
  wire [31:0] R7269;
  wire [31:0] R7268;
  wire [31:0] R7267;
  wire [31:0] R7266;
  wire [31:0] R7265;
  wire [31:0] R7264;
  wire [31:0] R7263;
  wire [31:0] R7262;
  wire [31:0] R7261;
  wire [31:0] R7260;
  wire [31:0] R7259;
  wire [31:0] R7258;
  wire [31:0] R7257;
  wire [31:0] R7256;
  wire [31:0] R7255;
  wire [31:0] R7254;
  wire [31:0] R7253;
  wire [31:0] R7252;
  wire [31:0] R7251;
  wire [31:0] R7250;
  wire [31:0] R7249;
  wire [31:0] R7248;
  wire [31:0] R7247;
  wire [31:0] R7246;
  wire [31:0] R7245;
  wire [31:0] R7244;
  wire [31:0] R7243;
  wire [31:0] R7242;
  wire [31:0] R7241;
  wire [31:0] R7240;
  wire [31:0] R7239;
  wire [31:0] R7238;
  wire [31:0] R7237;
  wire [31:0] R7236;
  wire [31:0] R7235;
  wire [31:0] R7234;
  wire [31:0] R7233;
  wire [31:0] R7232;
  wire [31:0] R7231;
  wire [31:0] R7230;
  wire [31:0] R7229;
  wire [31:0] R7228;
  wire [31:0] R7227;
  wire [31:0] R7226;
  wire [31:0] R7225;
  wire [31:0] R7224;
  wire [31:0] R7223;
  wire [31:0] R7222;
  wire [31:0] R7221;
  wire [31:0] R7220;
  wire [31:0] R7219;
  wire [31:0] R7218;
  wire [31:0] R7217;
  wire [31:0] R7216;
  wire [31:0] R7215;
  wire [31:0] R7214;
  wire [31:0] R7213;
  wire [31:0] R7212;
  wire [31:0] R7211;
  wire [31:0] R7210;
  wire [31:0] R7209;
  wire [31:0] R7208;
  wire [31:0] R7207;
  wire [31:0] R7206;
  wire [31:0] R7205;
  wire [31:0] R7204;
  wire [31:0] R7203;
  wire [31:0] R7202;
  wire [31:0] R7201;
  wire [31:0] R7200;
  wire [31:0] R7199;
  wire [31:0] R7198;
  wire [31:0] R7197;
  wire [31:0] R7196;
  wire [31:0] R7195;
  wire [31:0] R7194;
  wire [31:0] R7193;
  wire [31:0] R7192;
  wire [31:0] R7191;
  wire [31:0] R7190;
  wire [31:0] R7189;
  wire [31:0] R7188;
  wire [31:0] R7187;
  wire [31:0] R7186;
  wire [31:0] R7185;
  wire [31:0] R7184;
  wire [31:0] R7183;
  wire [31:0] R7182;
  wire [31:0] R7181;
  wire [31:0] R7180;
  wire [31:0] R7179;
  wire [31:0] R7178;
  wire [31:0] R7177;
  wire [31:0] R7176;
  wire [31:0] R7175;
  wire [31:0] R7174;
  wire [31:0] R7173;
  wire [31:0] R7172;
  wire [31:0] R7171;
  wire [31:0] R7170;
  wire [31:0] R7169;
  wire [31:0] R7168;
  wire [31:0] R7167;
  wire [31:0] R7166;
  wire [31:0] R7165;
  wire [31:0] R7164;
  wire [31:0] R7163;
  wire [31:0] R7162;
  wire [31:0] R7161;
  wire [31:0] R7160;
  wire [31:0] R7159;
  wire [31:0] R7158;
  wire [31:0] R7157;
  wire [31:0] R7156;
  wire [31:0] R7155;
  wire [31:0] R7154;
  wire [31:0] R7153;
  wire [31:0] R7152;
  wire [31:0] R7151;
  wire [31:0] R7150;
  wire [31:0] R7149;
  wire [31:0] R7148;
  wire [31:0] R7147;
  wire [31:0] R7146;
  wire [31:0] R7145;
  wire [31:0] R7144;
  wire [31:0] R7143;
  wire [31:0] R7142;
  wire [31:0] R7141;
  wire [31:0] R7140;
  wire [31:0] R7139;
  wire [31:0] R7138;
  wire [31:0] R7137;
  wire [31:0] R7136;
  wire [31:0] R7135;
  wire [31:0] R7134;
  wire [31:0] R7133;
  wire [31:0] R7132;
  wire [31:0] R7131;
  wire [31:0] R7130;
  wire [31:0] R7129;
  wire [31:0] R7128;
  wire [31:0] R7127;
  wire [31:0] R7126;
  wire [31:0] R7125;
  wire [31:0] R7124;
  wire [31:0] R7123;
  wire [31:0] R7122;
  wire [31:0] R7121;
  wire [31:0] R7120;
  wire [31:0] R7119;
  wire [31:0] R7118;
  wire [31:0] R7117;
  wire [31:0] R7116;
  wire [31:0] R7115;
  wire [31:0] R7114;
  wire [31:0] R7113;
  wire [31:0] R7112;
  wire [31:0] R7111;
  wire [31:0] R7110;
  wire [31:0] R7109;
  wire [31:0] R7108;
  wire [31:0] R7107;
  wire [31:0] R7106;
  wire [31:0] R7105;
  wire [31:0] R7104;
  wire [31:0] R7103;
  wire [63:0] R7102;
  wire [31:0] R7101;
  wire [63:0] R7100;
  wire [63:0] R7099;
  wire [63:0] R7098;
  wire [63:0] R7097;
  wire [63:0] R7096;
  wire [63:0] R7095;
  wire [63:0] R7094;
  wire [63:0] R7093;
  wire [63:0] R7092;
  wire [63:0] R7091;
  wire [63:0] R7090;
  wire [63:0] R7089;
  wire [63:0] R7088;
  wire [63:0] R7087;
  wire [63:0] R7086;
  wire [63:0] R7085;
  wire [63:0] R7084;
  wire [63:0] R7083;
  wire [63:0] R7082;
  wire [63:0] R7081;
  wire [63:0] R7080;
  wire [63:0] R7079;
  wire [63:0] R7078;
  wire [63:0] R7077;
  wire [63:0] R7076;
  wire [63:0] R7075;
  wire [63:0] R7074;
  wire [63:0] R7073;
  wire [63:0] R7072;
  wire [63:0] R7071;
  wire [63:0] R7070;
  wire [63:0] R7069;
  wire [63:0] R7068;
  wire [63:0] R7067;
  wire [63:0] R7066;
  wire [63:0] R7065;
  wire [63:0] R7064;
  wire [63:0] R7063;
  wire [63:0] R7062;
  wire [63:0] R7061;
  wire [63:0] R7060;
  wire [63:0] R7059;
  wire [63:0] R7058;
  wire [63:0] R7057;
  wire [63:0] R7056;
  wire [63:0] R7055;
  wire [0:0] R7054;
  wire [0:0] R7053;
  wire [0:0] R7052;
  wire [0:0] R7051;
  wire [0:0] R7050;
  wire [0:0] R7049;
  wire [0:0] R7048;
  wire [0:0] R7047;
  wire [0:0] R7046;
  wire [0:0] R7045;
  wire [0:0] R7044;
  wire [0:0] R7043;
  wire [0:0] R7042;
  wire [0:0] R7041;
  wire [0:0] R7040;
  wire [0:0] R7039;
  wire [0:0] R7038;
  wire [0:0] R7037;
  wire [0:0] R7036;
  wire [0:0] R7035;
  wire [0:0] R7034;
  wire [0:0] R7033;
  wire [0:0] R7032;
  wire [0:0] R7031;
  wire [0:0] R7030;
  wire [0:0] R7029;
  wire [0:0] R7028;
  wire [0:0] R7027;
  wire [0:0] R7026;
  wire [0:0] R7025;
  wire [0:0] R7024;
  wire [0:0] R7023;
  wire [0:0] R7022;
  wire [0:0] R7021;
  wire [0:0] R7020;
  wire [0:0] R7019;
  wire [0:0] R7018;
  wire [0:0] R7017;
  wire [0:0] R7016;
  wire [0:0] R7015;
  wire [0:0] R7014;
  wire [0:0] R7013;
  wire [0:0] R7012;
  wire [0:0] R7011;
  wire [0:0] R7010;
  wire [0:0] R7009;
  wire [0:0] R7008;
  wire [0:0] R7007;
  wire [0:0] R7006;
  wire [0:0] R7005;
  wire [0:0] R7004;
  wire [0:0] R7003;
  wire [0:0] R7002;
  wire [0:0] R7001;
  wire [0:0] R7000;
  wire [0:0] R6999;
  wire [0:0] R6998;
  wire [0:0] R6997;
  wire [0:0] R6996;
  wire [0:0] R6995;
  wire [0:0] R6994;
  wire [0:0] R6993;
  wire [0:0] R6992;
  wire [0:0] R6991;
  wire [0:0] R6990;
  wire [0:0] R6989;
  wire [0:0] R6988;
  wire [0:0] R6987;
  wire [0:0] R6986;
  wire [0:0] R6985;
  wire [0:0] R6984;
  wire [0:0] R6983;
  wire [0:0] R6982;
  wire [0:0] R6981;
  wire [0:0] R6980;
  wire [0:0] R6979;
  wire [0:0] R6978;
  wire [0:0] R6977;
  wire [0:0] R6976;
  wire [0:0] R6975;
  wire [0:0] R6974;
  wire [0:0] R6973;
  wire [0:0] R6972;
  wire [0:0] R6971;
  wire [0:0] R6970;
  wire [0:0] R6969;
  wire [0:0] R6968;
  wire [0:0] R6967;
  wire [0:0] R6966;
  wire [0:0] R6965;
  wire [0:0] R6964;
  wire [0:0] R6963;
  wire [0:0] R6962;
  wire [0:0] R6961;
  wire [0:0] R6960;
  wire [0:0] R6959;
  wire [0:0] R6958;
  wire [0:0] R6957;
  wire [0:0] R6956;
  wire [0:0] R6955;
  wire [0:0] R6954;
  wire [0:0] R6953;
  wire [0:0] R6952;
  wire [0:0] R6951;
  wire [0:0] R6950;
  wire [0:0] R6949;
  wire [0:0] R6948;
  wire [0:0] R6947;
  wire [0:0] R6946;
  wire [0:0] R6945;
  wire [0:0] R6944;
  wire [0:0] R6943;
  wire [0:0] R6942;
  wire [0:0] R6941;
  wire [0:0] R6940;
  wire [0:0] R6939;
  wire [0:0] R6938;
  wire [0:0] R6937;
  wire [0:0] R6936;
  wire [0:0] R6935;
  wire [0:0] R6934;
  wire [0:0] R6933;
  wire [0:0] R6932;
  wire [0:0] R6931;
  wire [0:0] R6930;
  wire [0:0] R6929;
  wire [0:0] R6928;
  wire [0:0] R6927;
  wire [0:0] R6926;
  wire [0:0] R6925;
  wire [0:0] R6924;
  wire [0:0] R6923;
  wire [0:0] R6922;
  wire [0:0] R6921;
  wire [0:0] R6920;
  wire [0:0] R6919;
  wire [0:0] R6918;
  wire [0:0] R6917;
  wire [0:0] R6916;
  wire [0:0] R6915;
  wire [0:0] R6914;
  wire [0:0] R6913;
  wire [0:0] R6912;
  wire [0:0] R6911;
  wire [0:0] R6910;
  wire [0:0] R6909;
  wire [0:0] R6908;
  wire [0:0] R6907;
  wire [0:0] R6906;
  wire [0:0] R6905;
  wire [0:0] R6904;
  wire [0:0] R6903;
  wire [0:0] R6902;
  wire [0:0] R6901;
  wire [0:0] R6900;
  wire [0:0] R6899;
  wire [0:0] R6898;
  wire [0:0] R6897;
  wire [0:0] R6896;
  wire [0:0] R6895;
  wire [0:0] R6894;
  wire [0:0] R6893;
  wire [0:0] R6892;
  wire [0:0] R6891;
  wire [0:0] R6890;
  wire [0:0] R6889;
  wire [0:0] R6888;
  wire [0:0] R6887;
  wire [0:0] R6886;
  wire [0:0] R6885;
  wire [0:0] R6884;
  wire [0:0] R6883;
  wire [0:0] R6882;
  wire [0:0] R6881;
  wire [0:0] R6880;
  wire [0:0] R6879;
  wire [0:0] R6878;
  wire [0:0] R6877;
  wire [0:0] R6876;
  wire [0:0] R6875;
  wire [0:0] R6874;
  wire [0:0] R6873;
  wire [0:0] R6872;
  wire [0:0] R6871;
  wire [0:0] R6870;
  wire [0:0] R6869;
  wire [0:0] R6868;
  wire [0:0] R6867;
  wire [0:0] R6866;
  wire [0:0] R6865;
  wire [0:0] R6864;
  wire [0:0] R6863;
  wire [0:0] R6862;
  wire [0:0] R6861;
  wire [0:0] R6860;
  wire [0:0] R6859;
  wire [0:0] R6858;
  wire [0:0] R6857;
  wire [0:0] R6856;
  wire [0:0] R6855;
  wire [0:0] R6854;
  wire [0:0] R6853;
  wire [0:0] R6852;
  wire [0:0] R6851;
  wire [0:0] R6850;
  wire [0:0] R6849;
  wire [0:0] R6848;
  wire [63:0] R6847;
  wire [31:0] R6846;
  wire [31:0] R6845;
  wire [31:0] R6844;
  wire [31:0] R6843;
  wire [31:0] R6842;
  wire [31:0] R6841;
  wire [31:0] R6840;
  wire [31:0] R6839;
  wire [31:0] R6838;
  wire [31:0] R6837;
  wire [31:0] R6836;
  wire [31:0] R6835;
  wire [31:0] R6834;
  wire [31:0] R6833;
  wire [31:0] R6832;
  wire [31:0] R6831;
  wire [31:0] R6830;
  wire [31:0] R6829;
  wire [31:0] R6828;
  wire [31:0] R6827;
  wire [31:0] R6826;
  wire [31:0] R6825;
  wire [31:0] R6824;
  wire [31:0] R6823;
  wire [31:0] R6822;
  wire [31:0] R6821;
  wire [31:0] R6820;
  wire [31:0] R6819;
  wire [31:0] R6818;
  wire [31:0] R6817;
  wire [31:0] R6816;
  wire [31:0] R6815;
  wire [31:0] R6814;
  wire [31:0] R6813;
  wire [31:0] R6812;
  wire [31:0] R6811;
  wire [31:0] R6810;
  wire [31:0] R6809;
  wire [31:0] R6808;
  wire [31:0] R6807;
  wire [31:0] R6806;
  wire [31:0] R6805;
  wire [31:0] R6804;
  wire [31:0] R6803;
  wire [31:0] R6802;
  wire [31:0] R6801;
  wire [31:0] R6800;
  wire [31:0] R6799;
  wire [31:0] R6798;
  wire [31:0] R6797;
  wire [31:0] R6796;
  wire [31:0] R6795;
  wire [31:0] R6794;
  wire [31:0] R6793;
  wire [31:0] R6792;
  wire [31:0] R6791;
  wire [31:0] R6790;
  wire [31:0] R6789;
  wire [31:0] R6788;
  wire [31:0] R6787;
  wire [31:0] R6786;
  wire [31:0] R6785;
  wire [31:0] R6784;
  wire [31:0] R6783;
  wire [31:0] R6782;
  wire [31:0] R6781;
  wire [31:0] R6780;
  wire [31:0] R6779;
  wire [31:0] R6778;
  wire [31:0] R6777;
  wire [31:0] R6776;
  wire [31:0] R6775;
  wire [31:0] R6774;
  wire [31:0] R6773;
  wire [31:0] R6772;
  wire [31:0] R6771;
  wire [31:0] R6770;
  wire [31:0] R6769;
  wire [31:0] R6768;
  wire [31:0] R6767;
  wire [31:0] R6766;
  wire [31:0] R6765;
  wire [31:0] R6764;
  wire [31:0] R6763;
  wire [31:0] R6762;
  wire [31:0] R6761;
  wire [31:0] R6760;
  wire [31:0] R6759;
  wire [31:0] R6758;
  wire [31:0] R6757;
  wire [31:0] R6756;
  wire [31:0] R6755;
  wire [31:0] R6754;
  wire [31:0] R6753;
  wire [31:0] R6752;
  wire [31:0] R6751;
  wire [31:0] R6750;
  wire [31:0] R6749;
  wire [31:0] R6748;
  wire [31:0] R6747;
  wire [31:0] R6746;
  wire [31:0] R6745;
  wire [31:0] R6744;
  wire [31:0] R6743;
  wire [31:0] R6742;
  wire [31:0] R6741;
  wire [31:0] R6740;
  wire [31:0] R6739;
  wire [31:0] R6738;
  wire [31:0] R6737;
  wire [31:0] R6736;
  wire [31:0] R6735;
  wire [31:0] R6734;
  wire [31:0] R6733;
  wire [31:0] R6732;
  wire [31:0] R6731;
  wire [31:0] R6730;
  wire [31:0] R6729;
  wire [31:0] R6728;
  wire [31:0] R6727;
  wire [31:0] R6726;
  wire [31:0] R6725;
  wire [31:0] R6724;
  wire [31:0] R6723;
  wire [31:0] R6722;
  wire [31:0] R6721;
  wire [31:0] R6720;
  wire [31:0] R6719;
  wire [31:0] R6718;
  wire [31:0] R6717;
  wire [31:0] R6716;
  wire [31:0] R6715;
  wire [31:0] R6714;
  wire [31:0] R6713;
  wire [31:0] R6712;
  wire [31:0] R6711;
  wire [31:0] R6710;
  wire [31:0] R6709;
  wire [31:0] R6708;
  wire [31:0] R6707;
  wire [31:0] R6706;
  wire [31:0] R6705;
  wire [31:0] R6704;
  wire [31:0] R6703;
  wire [31:0] R6702;
  wire [31:0] R6701;
  wire [31:0] R6700;
  wire [31:0] R6699;
  wire [31:0] R6698;
  wire [31:0] R6697;
  wire [31:0] R6696;
  wire [31:0] R6695;
  wire [31:0] R6694;
  wire [31:0] R6693;
  wire [31:0] R6692;
  wire [31:0] R6691;
  wire [31:0] R6690;
  wire [31:0] R6689;
  wire [31:0] R6688;
  wire [31:0] R6687;
  wire [31:0] R6686;
  wire [31:0] R6685;
  wire [31:0] R6684;
  wire [31:0] R6683;
  wire [31:0] R6682;
  wire [31:0] R6681;
  wire [31:0] R6680;
  wire [31:0] R6679;
  wire [31:0] R6678;
  wire [31:0] R6677;
  wire [31:0] R6676;
  wire [31:0] R6675;
  wire [31:0] R6674;
  wire [31:0] R6673;
  wire [31:0] R6672;
  wire [31:0] R6671;
  wire [31:0] R6670;
  wire [31:0] R6669;
  wire [31:0] R6668;
  wire [31:0] R6667;
  wire [31:0] R6666;
  wire [31:0] R6665;
  wire [31:0] R6664;
  wire [31:0] R6663;
  wire [31:0] R6662;
  wire [31:0] R6661;
  wire [31:0] R6660;
  wire [31:0] R6659;
  wire [31:0] R6658;
  wire [31:0] R6657;
  wire [31:0] R6656;
  wire [31:0] R6655;
  wire [31:0] R6654;
  wire [31:0] R6653;
  wire [31:0] R6652;
  wire [31:0] R6651;
  wire [31:0] R6650;
  wire [31:0] R6649;
  wire [31:0] R6648;
  wire [31:0] R6647;
  wire [63:0] R6646;
  wire [63:0] R6645;
  wire [63:0] R6644;
  wire [31:0] R6643;
  wire [31:0] R6642;
  wire [31:0] R6641;
  wire [31:0] R6640;
  wire [31:0] R6639;
  wire [31:0] R6638;
  wire [31:0] R6637;
  wire [31:0] R6636;
  wire [31:0] R6635;
  wire [31:0] R6634;
  wire [31:0] R6633;
  wire [31:0] R6632;
  wire [31:0] R6631;
  wire [31:0] R6630;
  wire [31:0] R6629;
  wire [31:0] R6628;
  wire [31:0] R6627;
  wire [31:0] R6626;
  wire [31:0] R6625;
  wire [31:0] R6624;
  wire [31:0] R6623;
  wire [31:0] R6622;
  wire [31:0] R6621;
  wire [31:0] R6620;
  wire [31:0] R6619;
  wire [31:0] R6618;
  wire [31:0] R6617;
  wire [31:0] R6616;
  wire [31:0] R6615;
  wire [31:0] R6614;
  wire [31:0] R6613;
  wire [31:0] R6612;
  wire [31:0] R6611;
  wire [31:0] R6610;
  wire [31:0] R6609;
  wire [31:0] R6608;
  wire [31:0] R6607;
  wire [31:0] R6606;
  wire [31:0] R6605;
  wire [31:0] R6604;
  wire [31:0] R6603;
  wire [31:0] R6602;
  wire [31:0] R6601;
  wire [31:0] R6600;
  wire [31:0] R6599;
  wire [31:0] R6598;
  wire [31:0] R6597;
  wire [31:0] R6596;
  wire [31:0] R6595;
  wire [31:0] R6594;
  wire [31:0] R6593;
  wire [31:0] R6592;
  wire [31:0] R6591;
  wire [31:0] R6590;
  wire [31:0] R6589;
  wire [31:0] R6588;
  wire [31:0] R6587;
  wire [31:0] R6586;
  wire [31:0] R6585;
  wire [31:0] R6584;
  wire [31:0] R6583;
  wire [31:0] R6582;
  wire [31:0] R6581;
  wire [31:0] R6580;
  wire [31:0] R6579;
  wire [31:0] R6578;
  wire [31:0] R6577;
  wire [31:0] R6576;
  wire [31:0] R6575;
  wire [31:0] R6574;
  wire [31:0] R6573;
  wire [31:0] R6572;
  wire [31:0] R6571;
  wire [31:0] R6570;
  wire [31:0] R6569;
  wire [31:0] R6568;
  wire [31:0] R6567;
  wire [31:0] R6566;
  wire [31:0] R6565;
  wire [31:0] R6564;
  wire [31:0] R6563;
  wire [31:0] R6562;
  wire [31:0] R6561;
  wire [31:0] R6560;
  wire [31:0] R6559;
  wire [31:0] R6558;
  wire [31:0] R6557;
  wire [31:0] R6556;
  wire [31:0] R6555;
  wire [31:0] R6554;
  wire [31:0] R6553;
  wire [31:0] R6552;
  wire [31:0] R6551;
  wire [31:0] R6550;
  wire [31:0] R6549;
  wire [31:0] R6548;
  wire [31:0] R6547;
  wire [31:0] R6546;
  wire [31:0] R6545;
  wire [31:0] R6544;
  wire [31:0] R6543;
  wire [31:0] R6542;
  wire [31:0] R6541;
  wire [31:0] R6540;
  wire [31:0] R6539;
  wire [31:0] R6538;
  wire [31:0] R6537;
  wire [31:0] R6536;
  wire [31:0] R6535;
  wire [31:0] R6534;
  wire [31:0] R6533;
  wire [31:0] R6532;
  wire [31:0] R6531;
  wire [31:0] R6530;
  wire [31:0] R6529;
  wire [31:0] R6528;
  wire [31:0] R6527;
  wire [31:0] R6526;
  wire [31:0] R6525;
  wire [31:0] R6524;
  wire [31:0] R6523;
  wire [31:0] R6522;
  wire [31:0] R6521;
  wire [31:0] R6520;
  wire [31:0] R6519;
  wire [31:0] R6518;
  wire [31:0] R6517;
  wire [31:0] R6516;
  wire [31:0] R6515;
  wire [31:0] R6514;
  wire [31:0] R6513;
  wire [31:0] R6512;
  wire [31:0] R6511;
  wire [31:0] R6510;
  wire [31:0] R6509;
  wire [31:0] R6508;
  wire [31:0] R6507;
  wire [31:0] R6506;
  wire [31:0] R6505;
  wire [31:0] R6504;
  wire [31:0] R6503;
  wire [31:0] R6502;
  wire [31:0] R6501;
  wire [31:0] R6500;
  wire [31:0] R6499;
  wire [31:0] R6498;
  wire [31:0] R6497;
  wire [31:0] R6496;
  wire [31:0] R6495;
  wire [31:0] R6494;
  wire [31:0] R6493;
  wire [31:0] R6492;
  wire [31:0] R6491;
  wire [31:0] R6490;
  wire [31:0] R6489;
  wire [31:0] R6488;
  wire [31:0] R6487;
  wire [31:0] R6486;
  wire [31:0] R6485;
  wire [31:0] R6484;
  wire [31:0] R6483;
  wire [31:0] R6482;
  wire [31:0] R6481;
  wire [31:0] R6480;
  wire [31:0] R6479;
  wire [31:0] R6478;
  wire [31:0] R6477;
  wire [31:0] R6476;
  wire [31:0] R6475;
  wire [31:0] R6474;
  wire [31:0] R6473;
  wire [31:0] R6472;
  wire [31:0] R6471;
  wire [31:0] R6470;
  wire [31:0] R6469;
  wire [31:0] R6468;
  wire [31:0] R6467;
  wire [31:0] R6466;
  wire [31:0] R6465;
  wire [31:0] R6464;
  wire [31:0] R6463;
  wire [31:0] R6462;
  wire [31:0] R6461;
  wire [31:0] R6460;
  wire [31:0] R6459;
  wire [31:0] R6458;
  wire [31:0] R6457;
  wire [31:0] R6456;
  wire [31:0] R6455;
  wire [31:0] R6454;
  wire [31:0] R6453;
  wire [31:0] R6452;
  wire [31:0] R6451;
  wire [31:0] R6450;
  wire [31:0] R6449;
  wire [31:0] R6448;
  wire [31:0] R6447;
  wire [31:0] R6446;
  wire [31:0] R6445;
  wire [31:0] R6444;
  wire [31:0] R6443;
  wire [31:0] R6442;
  wire [31:0] R6441;
  wire [31:0] R6440;
  wire [31:0] R6439;
  wire [31:0] R6438;
  wire [63:0] R6437;
  wire [31:0] R6436;
  wire [63:0] R6435;
  wire [63:0] R6434;
  wire [63:0] R6433;
  wire [63:0] R6432;
  wire [63:0] R6431;
  wire [63:0] R6430;
  wire [63:0] R6429;
  wire [63:0] R6428;
  wire [63:0] R6427;
  wire [63:0] R6426;
  wire [63:0] R6425;
  wire [63:0] R6424;
  wire [63:0] R6423;
  wire [63:0] R6422;
  wire [63:0] R6421;
  wire [63:0] R6420;
  wire [63:0] R6419;
  wire [63:0] R6418;
  wire [63:0] R6417;
  wire [63:0] R6416;
  wire [63:0] R6415;
  wire [63:0] R6414;
  wire [63:0] R6413;
  wire [63:0] R6412;
  wire [63:0] R6411;
  wire [63:0] R6410;
  wire [63:0] R6409;
  wire [63:0] R6408;
  wire [63:0] R6407;
  wire [63:0] R6406;
  wire [63:0] R6405;
  wire [63:0] R6404;
  wire [63:0] R6403;
  wire [63:0] R6402;
  wire [63:0] R6401;
  wire [63:0] R6400;
  wire [63:0] R6399;
  wire [63:0] R6398;
  wire [63:0] R6397;
  wire [63:0] R6396;
  wire [63:0] R6395;
  wire [63:0] R6394;
  wire [63:0] R6393;
  wire [63:0] R6392;
  wire [63:0] R6391;
  wire [63:0] R6390;
  wire [0:0] R6389;
  wire [0:0] R6388;
  wire [0:0] R6387;
  wire [0:0] R6386;
  wire [0:0] R6385;
  wire [0:0] R6384;
  wire [0:0] R6383;
  wire [0:0] R6382;
  wire [0:0] R6381;
  wire [0:0] R6380;
  wire [0:0] R6379;
  wire [0:0] R6378;
  wire [0:0] R6377;
  wire [0:0] R6376;
  wire [0:0] R6375;
  wire [0:0] R6374;
  wire [0:0] R6373;
  wire [0:0] R6372;
  wire [0:0] R6371;
  wire [0:0] R6370;
  wire [0:0] R6369;
  wire [0:0] R6368;
  wire [0:0] R6367;
  wire [0:0] R6366;
  wire [0:0] R6365;
  wire [0:0] R6364;
  wire [0:0] R6363;
  wire [0:0] R6362;
  wire [0:0] R6361;
  wire [0:0] R6360;
  wire [0:0] R6359;
  wire [0:0] R6358;
  wire [0:0] R6357;
  wire [0:0] R6356;
  wire [0:0] R6355;
  wire [0:0] R6354;
  wire [0:0] R6353;
  wire [0:0] R6352;
  wire [0:0] R6351;
  wire [0:0] R6350;
  wire [0:0] R6349;
  wire [0:0] R6348;
  wire [0:0] R6347;
  wire [0:0] R6346;
  wire [0:0] R6345;
  wire [0:0] R6344;
  wire [0:0] R6343;
  wire [0:0] R6342;
  wire [0:0] R6341;
  wire [0:0] R6340;
  wire [0:0] R6339;
  wire [0:0] R6338;
  wire [0:0] R6337;
  wire [0:0] R6336;
  wire [0:0] R6335;
  wire [0:0] R6334;
  wire [0:0] R6333;
  wire [0:0] R6332;
  wire [0:0] R6331;
  wire [0:0] R6330;
  wire [0:0] R6329;
  wire [0:0] R6328;
  wire [0:0] R6327;
  wire [0:0] R6326;
  wire [0:0] R6325;
  wire [0:0] R6324;
  wire [0:0] R6323;
  wire [0:0] R6322;
  wire [0:0] R6321;
  wire [0:0] R6320;
  wire [0:0] R6319;
  wire [0:0] R6318;
  wire [0:0] R6317;
  wire [0:0] R6316;
  wire [0:0] R6315;
  wire [0:0] R6314;
  wire [0:0] R6313;
  wire [0:0] R6312;
  wire [0:0] R6311;
  wire [0:0] R6310;
  wire [0:0] R6309;
  wire [0:0] R6308;
  wire [0:0] R6307;
  wire [0:0] R6306;
  wire [0:0] R6305;
  wire [0:0] R6304;
  wire [0:0] R6303;
  wire [0:0] R6302;
  wire [0:0] R6301;
  wire [0:0] R6300;
  wire [0:0] R6299;
  wire [0:0] R6298;
  wire [0:0] R6297;
  wire [0:0] R6296;
  wire [0:0] R6295;
  wire [0:0] R6294;
  wire [0:0] R6293;
  wire [0:0] R6292;
  wire [0:0] R6291;
  wire [0:0] R6290;
  wire [0:0] R6289;
  wire [0:0] R6288;
  wire [0:0] R6287;
  wire [0:0] R6286;
  wire [0:0] R6285;
  wire [0:0] R6284;
  wire [0:0] R6283;
  wire [0:0] R6282;
  wire [0:0] R6281;
  wire [0:0] R6280;
  wire [0:0] R6279;
  wire [0:0] R6278;
  wire [0:0] R6277;
  wire [0:0] R6276;
  wire [0:0] R6275;
  wire [0:0] R6274;
  wire [0:0] R6273;
  wire [0:0] R6272;
  wire [0:0] R6271;
  wire [0:0] R6270;
  wire [0:0] R6269;
  wire [0:0] R6268;
  wire [0:0] R6267;
  wire [0:0] R6266;
  wire [0:0] R6265;
  wire [0:0] R6264;
  wire [0:0] R6263;
  wire [0:0] R6262;
  wire [0:0] R6261;
  wire [0:0] R6260;
  wire [0:0] R6259;
  wire [0:0] R6258;
  wire [0:0] R6257;
  wire [0:0] R6256;
  wire [0:0] R6255;
  wire [0:0] R6254;
  wire [0:0] R6253;
  wire [0:0] R6252;
  wire [0:0] R6251;
  wire [0:0] R6250;
  wire [0:0] R6249;
  wire [0:0] R6248;
  wire [0:0] R6247;
  wire [0:0] R6246;
  wire [0:0] R6245;
  wire [0:0] R6244;
  wire [0:0] R6243;
  wire [0:0] R6242;
  wire [0:0] R6241;
  wire [0:0] R6240;
  wire [0:0] R6239;
  wire [0:0] R6238;
  wire [0:0] R6237;
  wire [0:0] R6236;
  wire [0:0] R6235;
  wire [0:0] R6234;
  wire [0:0] R6233;
  wire [0:0] R6232;
  wire [0:0] R6231;
  wire [0:0] R6230;
  wire [0:0] R6229;
  wire [0:0] R6228;
  wire [0:0] R6227;
  wire [0:0] R6226;
  wire [0:0] R6225;
  wire [0:0] R6224;
  wire [0:0] R6223;
  wire [0:0] R6222;
  wire [0:0] R6221;
  wire [0:0] R6220;
  wire [0:0] R6219;
  wire [0:0] R6218;
  wire [0:0] R6217;
  wire [0:0] R6216;
  wire [0:0] R6215;
  wire [0:0] R6214;
  wire [0:0] R6213;
  wire [0:0] R6212;
  wire [0:0] R6211;
  wire [0:0] R6210;
  wire [0:0] R6209;
  wire [0:0] R6208;
  wire [0:0] R6207;
  wire [0:0] R6206;
  wire [0:0] R6205;
  wire [0:0] R6204;
  wire [0:0] R6203;
  wire [0:0] R6202;
  wire [0:0] R6201;
  wire [0:0] R6200;
  wire [0:0] R6199;
  wire [0:0] R6198;
  wire [0:0] R6197;
  wire [0:0] R6196;
  wire [0:0] R6195;
  wire [0:0] R6194;
  wire [0:0] R6193;
  wire [0:0] R6192;
  wire [0:0] R6191;
  wire [0:0] R6190;
  wire [0:0] R6189;
  wire [0:0] R6188;
  wire [0:0] R6187;
  wire [0:0] R6186;
  wire [0:0] R6185;
  wire [0:0] R6184;
  wire [0:0] R6183;
  wire [0:0] R6182;
  wire [0:0] R6181;
  wire [0:0] R6180;
  wire [0:0] R6179;
  wire [0:0] R6178;
  wire [0:0] R6177;
  wire [0:0] R6176;
  wire [0:0] R6175;
  wire [0:0] R6174;
  wire [0:0] R6173;
  wire [0:0] R6172;
  wire [0:0] R6171;
  wire [0:0] R6170;
  wire [0:0] R6169;
  wire [63:0] R6168;
  wire [31:0] R6167;
  wire [31:0] R6166;
  wire [31:0] R6165;
  wire [31:0] R6164;
  wire [31:0] R6163;
  wire [31:0] R6162;
  wire [31:0] R6161;
  wire [31:0] R6160;
  wire [31:0] R6159;
  wire [31:0] R6158;
  wire [31:0] R6157;
  wire [31:0] R6156;
  wire [31:0] R6155;
  wire [31:0] R6154;
  wire [31:0] R6153;
  wire [31:0] R6152;
  wire [31:0] R6151;
  wire [31:0] R6150;
  wire [31:0] R6149;
  wire [31:0] R6148;
  wire [31:0] R6147;
  wire [31:0] R6146;
  wire [31:0] R6145;
  wire [31:0] R6144;
  wire [31:0] R6143;
  wire [31:0] R6142;
  wire [31:0] R6141;
  wire [31:0] R6140;
  wire [31:0] R6139;
  wire [31:0] R6138;
  wire [31:0] R6137;
  wire [31:0] R6136;
  wire [31:0] R6135;
  wire [31:0] R6134;
  wire [31:0] R6133;
  wire [31:0] R6132;
  wire [31:0] R6131;
  wire [31:0] R6130;
  wire [31:0] R6129;
  wire [31:0] R6128;
  wire [31:0] R6127;
  wire [31:0] R6126;
  wire [31:0] R6125;
  wire [31:0] R6124;
  wire [31:0] R6123;
  wire [31:0] R6122;
  wire [31:0] R6121;
  wire [31:0] R6120;
  wire [31:0] R6119;
  wire [31:0] R6118;
  wire [31:0] R6117;
  wire [31:0] R6116;
  wire [31:0] R6115;
  wire [31:0] R6114;
  wire [31:0] R6113;
  wire [31:0] R6112;
  wire [31:0] R6111;
  wire [31:0] R6110;
  wire [31:0] R6109;
  wire [31:0] R6108;
  wire [31:0] R6107;
  wire [31:0] R6106;
  wire [31:0] R6105;
  wire [31:0] R6104;
  wire [31:0] R6103;
  wire [31:0] R6102;
  wire [31:0] R6101;
  wire [31:0] R6100;
  wire [31:0] R6099;
  wire [31:0] R6098;
  wire [31:0] R6097;
  wire [31:0] R6096;
  wire [31:0] R6095;
  wire [31:0] R6094;
  wire [31:0] R6093;
  wire [31:0] R6092;
  wire [31:0] R6091;
  wire [31:0] R6090;
  wire [31:0] R6089;
  wire [31:0] R6088;
  wire [31:0] R6087;
  wire [31:0] R6086;
  wire [31:0] R6085;
  wire [31:0] R6084;
  wire [31:0] R6083;
  wire [31:0] R6082;
  wire [31:0] R6081;
  wire [31:0] R6080;
  wire [31:0] R6079;
  wire [31:0] R6078;
  wire [31:0] R6077;
  wire [31:0] R6076;
  wire [31:0] R6075;
  wire [31:0] R6074;
  wire [31:0] R6073;
  wire [31:0] R6072;
  wire [31:0] R6071;
  wire [31:0] R6070;
  wire [31:0] R6069;
  wire [31:0] R6068;
  wire [31:0] R6067;
  wire [31:0] R6066;
  wire [31:0] R6065;
  wire [31:0] R6064;
  wire [31:0] R6063;
  wire [31:0] R6062;
  wire [31:0] R6061;
  wire [31:0] R6060;
  wire [31:0] R6059;
  wire [31:0] R6058;
  wire [31:0] R6057;
  wire [31:0] R6056;
  wire [31:0] R6055;
  wire [31:0] R6054;
  wire [31:0] R6053;
  wire [31:0] R6052;
  wire [31:0] R6051;
  wire [31:0] R6050;
  wire [31:0] R6049;
  wire [31:0] R6048;
  wire [31:0] R6047;
  wire [31:0] R6046;
  wire [31:0] R6045;
  wire [31:0] R6044;
  wire [31:0] R6043;
  wire [31:0] R6042;
  wire [31:0] R6041;
  wire [31:0] R6040;
  wire [31:0] R6039;
  wire [31:0] R6038;
  wire [31:0] R6037;
  wire [31:0] R6036;
  wire [31:0] R6035;
  wire [31:0] R6034;
  wire [31:0] R6033;
  wire [31:0] R6032;
  wire [31:0] R6031;
  wire [31:0] R6030;
  wire [31:0] R6029;
  wire [31:0] R6028;
  wire [31:0] R6027;
  wire [31:0] R6026;
  wire [31:0] R6025;
  wire [31:0] R6024;
  wire [31:0] R6023;
  wire [31:0] R6022;
  wire [31:0] R6021;
  wire [31:0] R6020;
  wire [31:0] R6019;
  wire [31:0] R6018;
  wire [31:0] R6017;
  wire [31:0] R6016;
  wire [31:0] R6015;
  wire [31:0] R6014;
  wire [31:0] R6013;
  wire [31:0] R6012;
  wire [31:0] R6011;
  wire [31:0] R6010;
  wire [31:0] R6009;
  wire [31:0] R6008;
  wire [31:0] R6007;
  wire [31:0] R6006;
  wire [31:0] R6005;
  wire [31:0] R6004;
  wire [31:0] R6003;
  wire [31:0] R6002;
  wire [31:0] R6001;
  wire [31:0] R6000;
  wire [31:0] R5999;
  wire [31:0] R5998;
  wire [31:0] R5997;
  wire [31:0] R5996;
  wire [31:0] R5995;
  wire [31:0] R5994;
  wire [31:0] R5993;
  wire [31:0] R5992;
  wire [31:0] R5991;
  wire [31:0] R5990;
  wire [31:0] R5989;
  wire [31:0] R5988;
  wire [31:0] R5987;
  wire [31:0] R5986;
  wire [31:0] R5985;
  wire [31:0] R5984;
  wire [31:0] R5983;
  wire [31:0] R5982;
  wire [31:0] R5981;
  wire [31:0] R5980;
  wire [31:0] R5979;
  wire [31:0] R5978;
  wire [31:0] R5977;
  wire [31:0] R5976;
  wire [31:0] R5975;
  wire [31:0] R5974;
  wire [31:0] R5973;
  wire [31:0] R5972;
  wire [31:0] R5971;
  wire [31:0] R5970;
  wire [31:0] R5969;
  wire [31:0] R5968;
  wire [31:0] R5967;
  wire [31:0] R5966;
  wire [31:0] R5965;
  wire [31:0] R5964;
  wire [31:0] R5963;
  wire [31:0] R5962;
  wire [31:0] R5961;
  wire [31:0] R5960;
  wire [31:0] R5959;
  wire [31:0] R5958;
  wire [31:0] R5957;
  wire [31:0] R5956;
  wire [31:0] R5955;
  wire [63:0] R5954;
  wire [63:0] R5953;
  wire [63:0] R5952;
  wire [31:0] R5951;
  wire [31:0] R5950;
  wire [31:0] R5949;
  wire [31:0] R5948;
  wire [31:0] R5947;
  wire [31:0] R5946;
  wire [31:0] R5945;
  wire [31:0] R5944;
  wire [31:0] R5943;
  wire [31:0] R5942;
  wire [31:0] R5941;
  wire [31:0] R5940;
  wire [31:0] R5939;
  wire [31:0] R5938;
  wire [31:0] R5937;
  wire [31:0] R5936;
  wire [31:0] R5935;
  wire [31:0] R5934;
  wire [31:0] R5933;
  wire [31:0] R5932;
  wire [31:0] R5931;
  wire [31:0] R5930;
  wire [31:0] R5929;
  wire [31:0] R5928;
  wire [31:0] R5927;
  wire [31:0] R5926;
  wire [31:0] R5925;
  wire [31:0] R5924;
  wire [31:0] R5923;
  wire [31:0] R5922;
  wire [31:0] R5921;
  wire [31:0] R5920;
  wire [31:0] R5919;
  wire [31:0] R5918;
  wire [31:0] R5917;
  wire [31:0] R5916;
  wire [31:0] R5915;
  wire [31:0] R5914;
  wire [31:0] R5913;
  wire [31:0] R5912;
  wire [31:0] R5911;
  wire [31:0] R5910;
  wire [31:0] R5909;
  wire [31:0] R5908;
  wire [31:0] R5907;
  wire [31:0] R5906;
  wire [31:0] R5905;
  wire [31:0] R5904;
  wire [31:0] R5903;
  wire [31:0] R5902;
  wire [31:0] R5901;
  wire [31:0] R5900;
  wire [31:0] R5899;
  wire [31:0] R5898;
  wire [31:0] R5897;
  wire [31:0] R5896;
  wire [31:0] R5895;
  wire [31:0] R5894;
  wire [31:0] R5893;
  wire [31:0] R5892;
  wire [31:0] R5891;
  wire [31:0] R5890;
  wire [31:0] R5889;
  wire [31:0] R5888;
  wire [31:0] R5887;
  wire [31:0] R5886;
  wire [31:0] R5885;
  wire [31:0] R5884;
  wire [31:0] R5883;
  wire [31:0] R5882;
  wire [31:0] R5881;
  wire [31:0] R5880;
  wire [31:0] R5879;
  wire [31:0] R5878;
  wire [31:0] R5877;
  wire [31:0] R5876;
  wire [31:0] R5875;
  wire [31:0] R5874;
  wire [31:0] R5873;
  wire [31:0] R5872;
  wire [31:0] R5871;
  wire [31:0] R5870;
  wire [31:0] R5869;
  wire [31:0] R5868;
  wire [31:0] R5867;
  wire [31:0] R5866;
  wire [31:0] R5865;
  wire [31:0] R5864;
  wire [31:0] R5863;
  wire [31:0] R5862;
  wire [31:0] R5861;
  wire [31:0] R5860;
  wire [31:0] R5859;
  wire [31:0] R5858;
  wire [31:0] R5857;
  wire [31:0] R5856;
  wire [31:0] R5855;
  wire [31:0] R5854;
  wire [31:0] R5853;
  wire [31:0] R5852;
  wire [31:0] R5851;
  wire [31:0] R5850;
  wire [31:0] R5849;
  wire [31:0] R5848;
  wire [31:0] R5847;
  wire [31:0] R5846;
  wire [31:0] R5845;
  wire [31:0] R5844;
  wire [31:0] R5843;
  wire [31:0] R5842;
  wire [31:0] R5841;
  wire [31:0] R5840;
  wire [31:0] R5839;
  wire [31:0] R5838;
  wire [31:0] R5837;
  wire [31:0] R5836;
  wire [31:0] R5835;
  wire [31:0] R5834;
  wire [31:0] R5833;
  wire [31:0] R5832;
  wire [31:0] R5831;
  wire [31:0] R5830;
  wire [31:0] R5829;
  wire [31:0] R5828;
  wire [31:0] R5827;
  wire [31:0] R5826;
  wire [31:0] R5825;
  wire [31:0] R5824;
  wire [31:0] R5823;
  wire [31:0] R5822;
  wire [31:0] R5821;
  wire [31:0] R5820;
  wire [31:0] R5819;
  wire [31:0] R5818;
  wire [31:0] R5817;
  wire [31:0] R5816;
  wire [31:0] R5815;
  wire [31:0] R5814;
  wire [31:0] R5813;
  wire [31:0] R5812;
  wire [31:0] R5811;
  wire [31:0] R5810;
  wire [31:0] R5809;
  wire [31:0] R5808;
  wire [31:0] R5807;
  wire [31:0] R5806;
  wire [31:0] R5805;
  wire [31:0] R5804;
  wire [31:0] R5803;
  wire [31:0] R5802;
  wire [31:0] R5801;
  wire [31:0] R5800;
  wire [31:0] R5799;
  wire [31:0] R5798;
  wire [31:0] R5797;
  wire [31:0] R5796;
  wire [31:0] R5795;
  wire [31:0] R5794;
  wire [31:0] R5793;
  wire [31:0] R5792;
  wire [31:0] R5791;
  wire [31:0] R5790;
  wire [31:0] R5789;
  wire [31:0] R5788;
  wire [31:0] R5787;
  wire [31:0] R5786;
  wire [31:0] R5785;
  wire [31:0] R5784;
  wire [31:0] R5783;
  wire [31:0] R5782;
  wire [31:0] R5781;
  wire [31:0] R5780;
  wire [31:0] R5779;
  wire [31:0] R5778;
  wire [31:0] R5777;
  wire [31:0] R5776;
  wire [31:0] R5775;
  wire [31:0] R5774;
  wire [31:0] R5773;
  wire [31:0] R5772;
  wire [31:0] R5771;
  wire [31:0] R5770;
  wire [31:0] R5769;
  wire [31:0] R5768;
  wire [31:0] R5767;
  wire [31:0] R5766;
  wire [31:0] R5765;
  wire [31:0] R5764;
  wire [31:0] R5763;
  wire [31:0] R5762;
  wire [31:0] R5761;
  wire [31:0] R5760;
  wire [31:0] R5759;
  wire [31:0] R5758;
  wire [31:0] R5757;
  wire [31:0] R5756;
  wire [31:0] R5755;
  wire [31:0] R5754;
  wire [31:0] R5753;
  wire [31:0] R5752;
  wire [31:0] R5751;
  wire [31:0] R5750;
  wire [31:0] R5749;
  wire [31:0] R5748;
  wire [31:0] R5747;
  wire [31:0] R5746;
  wire [31:0] R5745;
  wire [31:0] R5744;
  wire [31:0] R5743;
  wire [31:0] R5742;
  wire [31:0] R5741;
  wire [31:0] R5740;
  wire [31:0] R5739;
  wire [31:0] R5738;
  wire [31:0] R5737;
  wire [31:0] R5736;
  wire [31:0] R5735;
  wire [31:0] R5734;
  wire [31:0] R5733;
  wire [63:0] R5732;
  wire [31:0] R5731;
  wire [63:0] R5730;
  wire [63:0] R5729;
  wire [63:0] R5728;
  wire [63:0] R5727;
  wire [63:0] R5726;
  wire [63:0] R5725;
  wire [63:0] R5724;
  wire [63:0] R5723;
  wire [63:0] R5722;
  wire [63:0] R5721;
  wire [63:0] R5720;
  wire [63:0] R5719;
  wire [63:0] R5718;
  wire [63:0] R5717;
  wire [63:0] R5716;
  wire [63:0] R5715;
  wire [63:0] R5714;
  wire [63:0] R5713;
  wire [63:0] R5712;
  wire [63:0] R5711;
  wire [63:0] R5710;
  wire [63:0] R5709;
  wire [63:0] R5708;
  wire [63:0] R5707;
  wire [63:0] R5706;
  wire [63:0] R5705;
  wire [63:0] R5704;
  wire [63:0] R5703;
  wire [63:0] R5702;
  wire [63:0] R5701;
  wire [63:0] R5700;
  wire [63:0] R5699;
  wire [63:0] R5698;
  wire [63:0] R5697;
  wire [63:0] R5696;
  wire [63:0] R5695;
  wire [63:0] R5694;
  wire [63:0] R5693;
  wire [63:0] R5692;
  wire [63:0] R5691;
  wire [63:0] R5690;
  wire [63:0] R5689;
  wire [63:0] R5688;
  wire [63:0] R5687;
  wire [63:0] R5686;
  wire [63:0] R5685;
  wire [0:0] R5684;
  wire [0:0] R5683;
  wire [0:0] R5682;
  wire [0:0] R5681;
  wire [0:0] R5680;
  wire [0:0] R5679;
  wire [0:0] R5678;
  wire [0:0] R5677;
  wire [0:0] R5676;
  wire [0:0] R5675;
  wire [0:0] R5674;
  wire [0:0] R5673;
  wire [0:0] R5672;
  wire [0:0] R5671;
  wire [0:0] R5670;
  wire [0:0] R5669;
  wire [0:0] R5668;
  wire [0:0] R5667;
  wire [0:0] R5666;
  wire [0:0] R5665;
  wire [0:0] R5664;
  wire [0:0] R5663;
  wire [0:0] R5662;
  wire [0:0] R5661;
  wire [0:0] R5660;
  wire [0:0] R5659;
  wire [0:0] R5658;
  wire [0:0] R5657;
  wire [0:0] R5656;
  wire [0:0] R5655;
  wire [0:0] R5654;
  wire [0:0] R5653;
  wire [0:0] R5652;
  wire [0:0] R5651;
  wire [0:0] R5650;
  wire [0:0] R5649;
  wire [0:0] R5648;
  wire [0:0] R5647;
  wire [0:0] R5646;
  wire [0:0] R5645;
  wire [0:0] R5644;
  wire [0:0] R5643;
  wire [0:0] R5642;
  wire [0:0] R5641;
  wire [0:0] R5640;
  wire [0:0] R5639;
  wire [0:0] R5638;
  wire [0:0] R5637;
  wire [0:0] R5636;
  wire [0:0] R5635;
  wire [0:0] R5634;
  wire [0:0] R5633;
  wire [0:0] R5632;
  wire [0:0] R5631;
  wire [0:0] R5630;
  wire [0:0] R5629;
  wire [0:0] R5628;
  wire [0:0] R5627;
  wire [0:0] R5626;
  wire [0:0] R5625;
  wire [0:0] R5624;
  wire [0:0] R5623;
  wire [0:0] R5622;
  wire [0:0] R5621;
  wire [0:0] R5620;
  wire [0:0] R5619;
  wire [0:0] R5618;
  wire [0:0] R5617;
  wire [0:0] R5616;
  wire [0:0] R5615;
  wire [0:0] R5614;
  wire [0:0] R5613;
  wire [0:0] R5612;
  wire [0:0] R5611;
  wire [0:0] R5610;
  wire [0:0] R5609;
  wire [0:0] R5608;
  wire [0:0] R5607;
  wire [0:0] R5606;
  wire [0:0] R5605;
  wire [0:0] R5604;
  wire [0:0] R5603;
  wire [0:0] R5602;
  wire [0:0] R5601;
  wire [0:0] R5600;
  wire [0:0] R5599;
  wire [0:0] R5598;
  wire [0:0] R5597;
  wire [0:0] R5596;
  wire [0:0] R5595;
  wire [0:0] R5594;
  wire [0:0] R5593;
  wire [0:0] R5592;
  wire [0:0] R5591;
  wire [0:0] R5590;
  wire [0:0] R5589;
  wire [0:0] R5588;
  wire [0:0] R5587;
  wire [0:0] R5586;
  wire [0:0] R5585;
  wire [0:0] R5584;
  wire [0:0] R5583;
  wire [0:0] R5582;
  wire [0:0] R5581;
  wire [0:0] R5580;
  wire [0:0] R5579;
  wire [0:0] R5578;
  wire [0:0] R5577;
  wire [0:0] R5576;
  wire [0:0] R5575;
  wire [0:0] R5574;
  wire [0:0] R5573;
  wire [0:0] R5572;
  wire [0:0] R5571;
  wire [0:0] R5570;
  wire [0:0] R5569;
  wire [0:0] R5568;
  wire [0:0] R5567;
  wire [0:0] R5566;
  wire [0:0] R5565;
  wire [0:0] R5564;
  wire [0:0] R5563;
  wire [0:0] R5562;
  wire [0:0] R5561;
  wire [0:0] R5560;
  wire [0:0] R5559;
  wire [0:0] R5558;
  wire [0:0] R5557;
  wire [0:0] R5556;
  wire [0:0] R5555;
  wire [0:0] R5554;
  wire [0:0] R5553;
  wire [0:0] R5552;
  wire [0:0] R5551;
  wire [0:0] R5550;
  wire [0:0] R5549;
  wire [0:0] R5548;
  wire [0:0] R5547;
  wire [0:0] R5546;
  wire [0:0] R5545;
  wire [0:0] R5544;
  wire [0:0] R5543;
  wire [0:0] R5542;
  wire [0:0] R5541;
  wire [0:0] R5540;
  wire [0:0] R5539;
  wire [0:0] R5538;
  wire [0:0] R5537;
  wire [0:0] R5536;
  wire [0:0] R5535;
  wire [0:0] R5534;
  wire [0:0] R5533;
  wire [0:0] R5532;
  wire [0:0] R5531;
  wire [0:0] R5530;
  wire [0:0] R5529;
  wire [0:0] R5528;
  wire [0:0] R5527;
  wire [0:0] R5526;
  wire [0:0] R5525;
  wire [0:0] R5524;
  wire [0:0] R5523;
  wire [0:0] R5522;
  wire [0:0] R5521;
  wire [0:0] R5520;
  wire [0:0] R5519;
  wire [0:0] R5518;
  wire [0:0] R5517;
  wire [0:0] R5516;
  wire [0:0] R5515;
  wire [0:0] R5514;
  wire [0:0] R5513;
  wire [0:0] R5512;
  wire [0:0] R5511;
  wire [0:0] R5510;
  wire [0:0] R5509;
  wire [0:0] R5508;
  wire [0:0] R5507;
  wire [0:0] R5506;
  wire [0:0] R5505;
  wire [0:0] R5504;
  wire [0:0] R5503;
  wire [0:0] R5502;
  wire [0:0] R5501;
  wire [0:0] R5500;
  wire [0:0] R5499;
  wire [0:0] R5498;
  wire [0:0] R5497;
  wire [0:0] R5496;
  wire [0:0] R5495;
  wire [0:0] R5494;
  wire [0:0] R5493;
  wire [0:0] R5492;
  wire [0:0] R5491;
  wire [0:0] R5490;
  wire [0:0] R5489;
  wire [0:0] R5488;
  wire [0:0] R5487;
  wire [0:0] R5486;
  wire [0:0] R5485;
  wire [0:0] R5484;
  wire [0:0] R5483;
  wire [0:0] R5482;
  wire [0:0] R5481;
  wire [0:0] R5480;
  wire [0:0] R5479;
  wire [0:0] R5478;
  wire [0:0] R5477;
  wire [0:0] R5476;
  wire [0:0] R5475;
  wire [0:0] R5474;
  wire [0:0] R5473;
  wire [0:0] R5472;
  wire [0:0] R5471;
  wire [0:0] R5470;
  wire [0:0] R5469;
  wire [0:0] R5468;
  wire [0:0] R5467;
  wire [0:0] R5466;
  wire [0:0] R5465;
  wire [0:0] R5464;
  wire [0:0] R5463;
  wire [0:0] R5462;
  wire [0:0] R5461;
  wire [0:0] R5460;
  wire [0:0] R5459;
  wire [0:0] R5458;
  wire [0:0] R5457;
  wire [0:0] R5456;
  wire [0:0] R5455;
  wire [0:0] R5454;
  wire [0:0] R5453;
  wire [0:0] R5452;
  wire [0:0] R5451;
  wire [63:0] R5450;
  wire [31:0] R5449;
  wire [31:0] R5448;
  wire [31:0] R5447;
  wire [31:0] R5446;
  wire [31:0] R5445;
  wire [31:0] R5444;
  wire [31:0] R5443;
  wire [31:0] R5442;
  wire [31:0] R5441;
  wire [31:0] R5440;
  wire [31:0] R5439;
  wire [31:0] R5438;
  wire [31:0] R5437;
  wire [31:0] R5436;
  wire [31:0] R5435;
  wire [31:0] R5434;
  wire [31:0] R5433;
  wire [31:0] R5432;
  wire [31:0] R5431;
  wire [31:0] R5430;
  wire [31:0] R5429;
  wire [31:0] R5428;
  wire [31:0] R5427;
  wire [31:0] R5426;
  wire [31:0] R5425;
  wire [31:0] R5424;
  wire [31:0] R5423;
  wire [31:0] R5422;
  wire [31:0] R5421;
  wire [31:0] R5420;
  wire [31:0] R5419;
  wire [31:0] R5418;
  wire [31:0] R5417;
  wire [31:0] R5416;
  wire [31:0] R5415;
  wire [31:0] R5414;
  wire [31:0] R5413;
  wire [31:0] R5412;
  wire [31:0] R5411;
  wire [31:0] R5410;
  wire [31:0] R5409;
  wire [31:0] R5408;
  wire [31:0] R5407;
  wire [31:0] R5406;
  wire [31:0] R5405;
  wire [31:0] R5404;
  wire [31:0] R5403;
  wire [31:0] R5402;
  wire [31:0] R5401;
  wire [31:0] R5400;
  wire [31:0] R5399;
  wire [31:0] R5398;
  wire [31:0] R5397;
  wire [31:0] R5396;
  wire [31:0] R5395;
  wire [31:0] R5394;
  wire [31:0] R5393;
  wire [31:0] R5392;
  wire [31:0] R5391;
  wire [31:0] R5390;
  wire [31:0] R5389;
  wire [31:0] R5388;
  wire [31:0] R5387;
  wire [31:0] R5386;
  wire [31:0] R5385;
  wire [31:0] R5384;
  wire [31:0] R5383;
  wire [31:0] R5382;
  wire [31:0] R5381;
  wire [31:0] R5380;
  wire [31:0] R5379;
  wire [31:0] R5378;
  wire [31:0] R5377;
  wire [31:0] R5376;
  wire [31:0] R5375;
  wire [31:0] R5374;
  wire [31:0] R5373;
  wire [31:0] R5372;
  wire [31:0] R5371;
  wire [31:0] R5370;
  wire [31:0] R5369;
  wire [31:0] R5368;
  wire [31:0] R5367;
  wire [31:0] R5366;
  wire [31:0] R5365;
  wire [31:0] R5364;
  wire [31:0] R5363;
  wire [31:0] R5362;
  wire [31:0] R5361;
  wire [31:0] R5360;
  wire [31:0] R5359;
  wire [31:0] R5358;
  wire [31:0] R5357;
  wire [31:0] R5356;
  wire [31:0] R5355;
  wire [31:0] R5354;
  wire [31:0] R5353;
  wire [31:0] R5352;
  wire [31:0] R5351;
  wire [31:0] R5350;
  wire [31:0] R5349;
  wire [31:0] R5348;
  wire [31:0] R5347;
  wire [31:0] R5346;
  wire [31:0] R5345;
  wire [31:0] R5344;
  wire [31:0] R5343;
  wire [31:0] R5342;
  wire [31:0] R5341;
  wire [31:0] R5340;
  wire [31:0] R5339;
  wire [31:0] R5338;
  wire [31:0] R5337;
  wire [31:0] R5336;
  wire [31:0] R5335;
  wire [31:0] R5334;
  wire [31:0] R5333;
  wire [31:0] R5332;
  wire [31:0] R5331;
  wire [31:0] R5330;
  wire [31:0] R5329;
  wire [31:0] R5328;
  wire [31:0] R5327;
  wire [31:0] R5326;
  wire [31:0] R5325;
  wire [31:0] R5324;
  wire [31:0] R5323;
  wire [31:0] R5322;
  wire [31:0] R5321;
  wire [31:0] R5320;
  wire [31:0] R5319;
  wire [31:0] R5318;
  wire [31:0] R5317;
  wire [31:0] R5316;
  wire [31:0] R5315;
  wire [31:0] R5314;
  wire [31:0] R5313;
  wire [31:0] R5312;
  wire [31:0] R5311;
  wire [31:0] R5310;
  wire [31:0] R5309;
  wire [31:0] R5308;
  wire [31:0] R5307;
  wire [31:0] R5306;
  wire [31:0] R5305;
  wire [31:0] R5304;
  wire [31:0] R5303;
  wire [31:0] R5302;
  wire [31:0] R5301;
  wire [31:0] R5300;
  wire [31:0] R5299;
  wire [31:0] R5298;
  wire [31:0] R5297;
  wire [31:0] R5296;
  wire [31:0] R5295;
  wire [31:0] R5294;
  wire [31:0] R5293;
  wire [31:0] R5292;
  wire [31:0] R5291;
  wire [31:0] R5290;
  wire [31:0] R5289;
  wire [31:0] R5288;
  wire [31:0] R5287;
  wire [31:0] R5286;
  wire [31:0] R5285;
  wire [31:0] R5284;
  wire [31:0] R5283;
  wire [31:0] R5282;
  wire [31:0] R5281;
  wire [31:0] R5280;
  wire [31:0] R5279;
  wire [31:0] R5278;
  wire [31:0] R5277;
  wire [31:0] R5276;
  wire [31:0] R5275;
  wire [31:0] R5274;
  wire [31:0] R5273;
  wire [31:0] R5272;
  wire [31:0] R5271;
  wire [31:0] R5270;
  wire [31:0] R5269;
  wire [31:0] R5268;
  wire [31:0] R5267;
  wire [31:0] R5266;
  wire [31:0] R5265;
  wire [31:0] R5264;
  wire [31:0] R5263;
  wire [31:0] R5262;
  wire [31:0] R5261;
  wire [31:0] R5260;
  wire [31:0] R5259;
  wire [31:0] R5258;
  wire [31:0] R5257;
  wire [31:0] R5256;
  wire [31:0] R5255;
  wire [31:0] R5254;
  wire [31:0] R5253;
  wire [31:0] R5252;
  wire [31:0] R5251;
  wire [31:0] R5250;
  wire [31:0] R5249;
  wire [31:0] R5248;
  wire [31:0] R5247;
  wire [31:0] R5246;
  wire [31:0] R5245;
  wire [31:0] R5244;
  wire [31:0] R5243;
  wire [31:0] R5242;
  wire [31:0] R5241;
  wire [31:0] R5240;
  wire [31:0] R5239;
  wire [31:0] R5238;
  wire [31:0] R5237;
  wire [31:0] R5236;
  wire [31:0] R5235;
  wire [31:0] R5234;
  wire [31:0] R5233;
  wire [31:0] R5232;
  wire [31:0] R5231;
  wire [31:0] R5230;
  wire [31:0] R5229;
  wire [31:0] R5228;
  wire [31:0] R5227;
  wire [31:0] R5226;
  wire [31:0] R5225;
  wire [31:0] R5224;
  wire [31:0] R5223;
  wire [63:0] R5222;
  wire [63:0] R5221;
  wire [63:0] R5220;
  wire [31:0] R5219;
  wire [31:0] R5218;
  wire [31:0] R5217;
  wire [31:0] R5216;
  wire [31:0] R5215;
  wire [31:0] R5214;
  wire [31:0] R5213;
  wire [31:0] R5212;
  wire [31:0] R5211;
  wire [31:0] R5210;
  wire [31:0] R5209;
  wire [31:0] R5208;
  wire [31:0] R5207;
  wire [31:0] R5206;
  wire [31:0] R5205;
  wire [31:0] R5204;
  wire [31:0] R5203;
  wire [31:0] R5202;
  wire [31:0] R5201;
  wire [31:0] R5200;
  wire [31:0] R5199;
  wire [31:0] R5198;
  wire [31:0] R5197;
  wire [31:0] R5196;
  wire [31:0] R5195;
  wire [31:0] R5194;
  wire [31:0] R5193;
  wire [31:0] R5192;
  wire [31:0] R5191;
  wire [31:0] R5190;
  wire [31:0] R5189;
  wire [31:0] R5188;
  wire [31:0] R5187;
  wire [31:0] R5186;
  wire [31:0] R5185;
  wire [31:0] R5184;
  wire [31:0] R5183;
  wire [31:0] R5182;
  wire [31:0] R5181;
  wire [31:0] R5180;
  wire [31:0] R5179;
  wire [31:0] R5178;
  wire [31:0] R5177;
  wire [31:0] R5176;
  wire [31:0] R5175;
  wire [31:0] R5174;
  wire [31:0] R5173;
  wire [31:0] R5172;
  wire [31:0] R5171;
  wire [31:0] R5170;
  wire [31:0] R5169;
  wire [31:0] R5168;
  wire [31:0] R5167;
  wire [31:0] R5166;
  wire [31:0] R5165;
  wire [31:0] R5164;
  wire [31:0] R5163;
  wire [31:0] R5162;
  wire [31:0] R5161;
  wire [31:0] R5160;
  wire [31:0] R5159;
  wire [31:0] R5158;
  wire [31:0] R5157;
  wire [31:0] R5156;
  wire [31:0] R5155;
  wire [31:0] R5154;
  wire [31:0] R5153;
  wire [31:0] R5152;
  wire [31:0] R5151;
  wire [31:0] R5150;
  wire [31:0] R5149;
  wire [31:0] R5148;
  wire [31:0] R5147;
  wire [31:0] R5146;
  wire [31:0] R5145;
  wire [31:0] R5144;
  wire [31:0] R5143;
  wire [31:0] R5142;
  wire [31:0] R5141;
  wire [31:0] R5140;
  wire [31:0] R5139;
  wire [31:0] R5138;
  wire [31:0] R5137;
  wire [31:0] R5136;
  wire [31:0] R5135;
  wire [31:0] R5134;
  wire [31:0] R5133;
  wire [31:0] R5132;
  wire [31:0] R5131;
  wire [31:0] R5130;
  wire [31:0] R5129;
  wire [31:0] R5128;
  wire [31:0] R5127;
  wire [31:0] R5126;
  wire [31:0] R5125;
  wire [31:0] R5124;
  wire [31:0] R5123;
  wire [31:0] R5122;
  wire [31:0] R5121;
  wire [31:0] R5120;
  wire [31:0] R5119;
  wire [31:0] R5118;
  wire [31:0] R5117;
  wire [31:0] R5116;
  wire [31:0] R5115;
  wire [31:0] R5114;
  wire [31:0] R5113;
  wire [31:0] R5112;
  wire [31:0] R5111;
  wire [31:0] R5110;
  wire [31:0] R5109;
  wire [31:0] R5108;
  wire [31:0] R5107;
  wire [31:0] R5106;
  wire [31:0] R5105;
  wire [31:0] R5104;
  wire [31:0] R5103;
  wire [31:0] R5102;
  wire [31:0] R5101;
  wire [31:0] R5100;
  wire [31:0] R5099;
  wire [31:0] R5098;
  wire [31:0] R5097;
  wire [31:0] R5096;
  wire [31:0] R5095;
  wire [31:0] R5094;
  wire [31:0] R5093;
  wire [31:0] R5092;
  wire [31:0] R5091;
  wire [31:0] R5090;
  wire [31:0] R5089;
  wire [31:0] R5088;
  wire [31:0] R5087;
  wire [31:0] R5086;
  wire [31:0] R5085;
  wire [31:0] R5084;
  wire [31:0] R5083;
  wire [31:0] R5082;
  wire [31:0] R5081;
  wire [31:0] R5080;
  wire [31:0] R5079;
  wire [31:0] R5078;
  wire [31:0] R5077;
  wire [31:0] R5076;
  wire [31:0] R5075;
  wire [31:0] R5074;
  wire [31:0] R5073;
  wire [31:0] R5072;
  wire [31:0] R5071;
  wire [31:0] R5070;
  wire [31:0] R5069;
  wire [31:0] R5068;
  wire [31:0] R5067;
  wire [31:0] R5066;
  wire [31:0] R5065;
  wire [31:0] R5064;
  wire [31:0] R5063;
  wire [31:0] R5062;
  wire [31:0] R5061;
  wire [31:0] R5060;
  wire [31:0] R5059;
  wire [31:0] R5058;
  wire [31:0] R5057;
  wire [31:0] R5056;
  wire [31:0] R5055;
  wire [31:0] R5054;
  wire [31:0] R5053;
  wire [31:0] R5052;
  wire [31:0] R5051;
  wire [31:0] R5050;
  wire [31:0] R5049;
  wire [31:0] R5048;
  wire [31:0] R5047;
  wire [31:0] R5046;
  wire [31:0] R5045;
  wire [31:0] R5044;
  wire [31:0] R5043;
  wire [31:0] R5042;
  wire [31:0] R5041;
  wire [31:0] R5040;
  wire [31:0] R5039;
  wire [31:0] R5038;
  wire [31:0] R5037;
  wire [31:0] R5036;
  wire [31:0] R5035;
  wire [31:0] R5034;
  wire [31:0] R5033;
  wire [31:0] R5032;
  wire [31:0] R5031;
  wire [31:0] R5030;
  wire [31:0] R5029;
  wire [31:0] R5028;
  wire [31:0] R5027;
  wire [31:0] R5026;
  wire [31:0] R5025;
  wire [31:0] R5024;
  wire [31:0] R5023;
  wire [31:0] R5022;
  wire [31:0] R5021;
  wire [31:0] R5020;
  wire [31:0] R5019;
  wire [31:0] R5018;
  wire [31:0] R5017;
  wire [31:0] R5016;
  wire [31:0] R5015;
  wire [31:0] R5014;
  wire [31:0] R5013;
  wire [31:0] R5012;
  wire [31:0] R5011;
  wire [31:0] R5010;
  wire [31:0] R5009;
  wire [31:0] R5008;
  wire [31:0] R5007;
  wire [31:0] R5006;
  wire [31:0] R5005;
  wire [31:0] R5004;
  wire [31:0] R5003;
  wire [31:0] R5002;
  wire [31:0] R5001;
  wire [31:0] R5000;
  wire [31:0] R4999;
  wire [31:0] R4998;
  wire [31:0] R4997;
  wire [31:0] R4996;
  wire [31:0] R4995;
  wire [31:0] R4994;
  wire [31:0] R4993;
  wire [31:0] R4992;
  wire [31:0] R4991;
  wire [31:0] R4990;
  wire [31:0] R4989;
  wire [31:0] R4988;
  wire [31:0] R4987;
  wire [63:0] R4986;
  wire [31:0] R4985;
  wire [63:0] R4984;
  wire [63:0] R4983;
  wire [63:0] R4982;
  wire [63:0] R4981;
  wire [63:0] R4980;
  wire [63:0] R4979;
  wire [63:0] R4978;
  wire [63:0] R4977;
  wire [63:0] R4976;
  wire [63:0] R4975;
  wire [63:0] R4974;
  wire [63:0] R4973;
  wire [63:0] R4972;
  wire [63:0] R4971;
  wire [63:0] R4970;
  wire [63:0] R4969;
  wire [63:0] R4968;
  wire [63:0] R4967;
  wire [63:0] R4966;
  wire [63:0] R4965;
  wire [63:0] R4964;
  wire [63:0] R4963;
  wire [63:0] R4962;
  wire [63:0] R4961;
  wire [63:0] R4960;
  wire [63:0] R4959;
  wire [63:0] R4958;
  wire [63:0] R4957;
  wire [63:0] R4956;
  wire [63:0] R4955;
  wire [63:0] R4954;
  wire [63:0] R4953;
  wire [63:0] R4952;
  wire [63:0] R4951;
  wire [63:0] R4950;
  wire [63:0] R4949;
  wire [63:0] R4948;
  wire [63:0] R4947;
  wire [63:0] R4946;
  wire [63:0] R4945;
  wire [63:0] R4944;
  wire [63:0] R4943;
  wire [63:0] R4942;
  wire [63:0] R4941;
  wire [63:0] R4940;
  wire [63:0] R4939;
  wire [0:0] R4938;
  wire [0:0] R4937;
  wire [0:0] R4936;
  wire [0:0] R4935;
  wire [0:0] R4934;
  wire [0:0] R4933;
  wire [0:0] R4932;
  wire [0:0] R4931;
  wire [0:0] R4930;
  wire [0:0] R4929;
  wire [0:0] R4928;
  wire [0:0] R4927;
  wire [0:0] R4926;
  wire [0:0] R4925;
  wire [0:0] R4924;
  wire [0:0] R4923;
  wire [0:0] R4922;
  wire [0:0] R4921;
  wire [0:0] R4920;
  wire [0:0] R4919;
  wire [0:0] R4918;
  wire [0:0] R4917;
  wire [0:0] R4916;
  wire [0:0] R4915;
  wire [0:0] R4914;
  wire [0:0] R4913;
  wire [0:0] R4912;
  wire [0:0] R4911;
  wire [0:0] R4910;
  wire [0:0] R4909;
  wire [0:0] R4908;
  wire [0:0] R4907;
  wire [0:0] R4906;
  wire [0:0] R4905;
  wire [0:0] R4904;
  wire [0:0] R4903;
  wire [0:0] R4902;
  wire [0:0] R4901;
  wire [0:0] R4900;
  wire [0:0] R4899;
  wire [0:0] R4898;
  wire [0:0] R4897;
  wire [0:0] R4896;
  wire [0:0] R4895;
  wire [0:0] R4894;
  wire [0:0] R4893;
  wire [0:0] R4892;
  wire [0:0] R4891;
  wire [0:0] R4890;
  wire [0:0] R4889;
  wire [0:0] R4888;
  wire [0:0] R4887;
  wire [0:0] R4886;
  wire [0:0] R4885;
  wire [0:0] R4884;
  wire [0:0] R4883;
  wire [0:0] R4882;
  wire [0:0] R4881;
  wire [0:0] R4880;
  wire [0:0] R4879;
  wire [0:0] R4878;
  wire [0:0] R4877;
  wire [0:0] R4876;
  wire [0:0] R4875;
  wire [0:0] R4874;
  wire [0:0] R4873;
  wire [0:0] R4872;
  wire [0:0] R4871;
  wire [0:0] R4870;
  wire [0:0] R4869;
  wire [0:0] R4868;
  wire [0:0] R4867;
  wire [0:0] R4866;
  wire [0:0] R4865;
  wire [0:0] R4864;
  wire [0:0] R4863;
  wire [0:0] R4862;
  wire [0:0] R4861;
  wire [0:0] R4860;
  wire [0:0] R4859;
  wire [0:0] R4858;
  wire [0:0] R4857;
  wire [0:0] R4856;
  wire [0:0] R4855;
  wire [0:0] R4854;
  wire [0:0] R4853;
  wire [0:0] R4852;
  wire [0:0] R4851;
  wire [0:0] R4850;
  wire [0:0] R4849;
  wire [0:0] R4848;
  wire [0:0] R4847;
  wire [0:0] R4846;
  wire [0:0] R4845;
  wire [0:0] R4844;
  wire [0:0] R4843;
  wire [0:0] R4842;
  wire [0:0] R4841;
  wire [0:0] R4840;
  wire [0:0] R4839;
  wire [0:0] R4838;
  wire [0:0] R4837;
  wire [0:0] R4836;
  wire [0:0] R4835;
  wire [0:0] R4834;
  wire [0:0] R4833;
  wire [0:0] R4832;
  wire [0:0] R4831;
  wire [0:0] R4830;
  wire [0:0] R4829;
  wire [0:0] R4828;
  wire [0:0] R4827;
  wire [0:0] R4826;
  wire [0:0] R4825;
  wire [0:0] R4824;
  wire [0:0] R4823;
  wire [0:0] R4822;
  wire [0:0] R4821;
  wire [0:0] R4820;
  wire [0:0] R4819;
  wire [0:0] R4818;
  wire [0:0] R4817;
  wire [0:0] R4816;
  wire [0:0] R4815;
  wire [0:0] R4814;
  wire [0:0] R4813;
  wire [0:0] R4812;
  wire [0:0] R4811;
  wire [0:0] R4810;
  wire [0:0] R4809;
  wire [0:0] R4808;
  wire [0:0] R4807;
  wire [0:0] R4806;
  wire [0:0] R4805;
  wire [0:0] R4804;
  wire [0:0] R4803;
  wire [0:0] R4802;
  wire [0:0] R4801;
  wire [0:0] R4800;
  wire [0:0] R4799;
  wire [0:0] R4798;
  wire [0:0] R4797;
  wire [0:0] R4796;
  wire [0:0] R4795;
  wire [0:0] R4794;
  wire [0:0] R4793;
  wire [0:0] R4792;
  wire [0:0] R4791;
  wire [0:0] R4790;
  wire [0:0] R4789;
  wire [0:0] R4788;
  wire [0:0] R4787;
  wire [0:0] R4786;
  wire [0:0] R4785;
  wire [0:0] R4784;
  wire [0:0] R4783;
  wire [0:0] R4782;
  wire [0:0] R4781;
  wire [0:0] R4780;
  wire [0:0] R4779;
  wire [0:0] R4778;
  wire [0:0] R4777;
  wire [0:0] R4776;
  wire [0:0] R4775;
  wire [0:0] R4774;
  wire [0:0] R4773;
  wire [0:0] R4772;
  wire [0:0] R4771;
  wire [0:0] R4770;
  wire [0:0] R4769;
  wire [0:0] R4768;
  wire [0:0] R4767;
  wire [0:0] R4766;
  wire [0:0] R4765;
  wire [0:0] R4764;
  wire [0:0] R4763;
  wire [0:0] R4762;
  wire [0:0] R4761;
  wire [0:0] R4760;
  wire [0:0] R4759;
  wire [0:0] R4758;
  wire [0:0] R4757;
  wire [0:0] R4756;
  wire [0:0] R4755;
  wire [0:0] R4754;
  wire [0:0] R4753;
  wire [0:0] R4752;
  wire [0:0] R4751;
  wire [0:0] R4750;
  wire [0:0] R4749;
  wire [0:0] R4748;
  wire [0:0] R4747;
  wire [0:0] R4746;
  wire [0:0] R4745;
  wire [0:0] R4744;
  wire [0:0] R4743;
  wire [0:0] R4742;
  wire [0:0] R4741;
  wire [0:0] R4740;
  wire [0:0] R4739;
  wire [0:0] R4738;
  wire [0:0] R4737;
  wire [0:0] R4736;
  wire [0:0] R4735;
  wire [0:0] R4734;
  wire [0:0] R4733;
  wire [0:0] R4732;
  wire [0:0] R4731;
  wire [0:0] R4730;
  wire [0:0] R4729;
  wire [0:0] R4728;
  wire [0:0] R4727;
  wire [0:0] R4726;
  wire [0:0] R4725;
  wire [0:0] R4724;
  wire [0:0] R4723;
  wire [0:0] R4722;
  wire [0:0] R4721;
  wire [0:0] R4720;
  wire [0:0] R4719;
  wire [0:0] R4718;
  wire [0:0] R4717;
  wire [0:0] R4716;
  wire [0:0] R4715;
  wire [0:0] R4714;
  wire [0:0] R4713;
  wire [0:0] R4712;
  wire [0:0] R4711;
  wire [0:0] R4710;
  wire [0:0] R4709;
  wire [0:0] R4708;
  wire [0:0] R4707;
  wire [0:0] R4706;
  wire [0:0] R4705;
  wire [0:0] R4704;
  wire [0:0] R4703;
  wire [0:0] R4702;
  wire [0:0] R4701;
  wire [0:0] R4700;
  wire [0:0] R4699;
  wire [0:0] R4698;
  wire [0:0] R4697;
  wire [0:0] R4696;
  wire [0:0] R4695;
  wire [0:0] R4694;
  wire [0:0] R4693;
  wire [0:0] R4692;
  wire [63:0] R4691;
  wire [31:0] R4690;
  wire [31:0] R4689;
  wire [31:0] R4688;
  wire [31:0] R4687;
  wire [31:0] R4686;
  wire [31:0] R4685;
  wire [31:0] R4684;
  wire [31:0] R4683;
  wire [31:0] R4682;
  wire [31:0] R4681;
  wire [31:0] R4680;
  wire [31:0] R4679;
  wire [31:0] R4678;
  wire [31:0] R4677;
  wire [31:0] R4676;
  wire [31:0] R4675;
  wire [31:0] R4674;
  wire [31:0] R4673;
  wire [31:0] R4672;
  wire [31:0] R4671;
  wire [31:0] R4670;
  wire [31:0] R4669;
  wire [31:0] R4668;
  wire [31:0] R4667;
  wire [31:0] R4666;
  wire [31:0] R4665;
  wire [31:0] R4664;
  wire [31:0] R4663;
  wire [31:0] R4662;
  wire [31:0] R4661;
  wire [31:0] R4660;
  wire [31:0] R4659;
  wire [31:0] R4658;
  wire [31:0] R4657;
  wire [31:0] R4656;
  wire [31:0] R4655;
  wire [31:0] R4654;
  wire [31:0] R4653;
  wire [31:0] R4652;
  wire [31:0] R4651;
  wire [31:0] R4650;
  wire [31:0] R4649;
  wire [31:0] R4648;
  wire [31:0] R4647;
  wire [31:0] R4646;
  wire [31:0] R4645;
  wire [31:0] R4644;
  wire [31:0] R4643;
  wire [31:0] R4642;
  wire [31:0] R4641;
  wire [31:0] R4640;
  wire [31:0] R4639;
  wire [31:0] R4638;
  wire [31:0] R4637;
  wire [31:0] R4636;
  wire [31:0] R4635;
  wire [31:0] R4634;
  wire [31:0] R4633;
  wire [31:0] R4632;
  wire [31:0] R4631;
  wire [31:0] R4630;
  wire [31:0] R4629;
  wire [31:0] R4628;
  wire [31:0] R4627;
  wire [31:0] R4626;
  wire [31:0] R4625;
  wire [31:0] R4624;
  wire [31:0] R4623;
  wire [31:0] R4622;
  wire [31:0] R4621;
  wire [31:0] R4620;
  wire [31:0] R4619;
  wire [31:0] R4618;
  wire [31:0] R4617;
  wire [31:0] R4616;
  wire [31:0] R4615;
  wire [31:0] R4614;
  wire [31:0] R4613;
  wire [31:0] R4612;
  wire [31:0] R4611;
  wire [31:0] R4610;
  wire [31:0] R4609;
  wire [31:0] R4608;
  wire [31:0] R4607;
  wire [31:0] R4606;
  wire [31:0] R4605;
  wire [31:0] R4604;
  wire [31:0] R4603;
  wire [31:0] R4602;
  wire [31:0] R4601;
  wire [31:0] R4600;
  wire [31:0] R4599;
  wire [31:0] R4598;
  wire [31:0] R4597;
  wire [31:0] R4596;
  wire [31:0] R4595;
  wire [31:0] R4594;
  wire [31:0] R4593;
  wire [31:0] R4592;
  wire [31:0] R4591;
  wire [31:0] R4590;
  wire [31:0] R4589;
  wire [31:0] R4588;
  wire [31:0] R4587;
  wire [31:0] R4586;
  wire [31:0] R4585;
  wire [31:0] R4584;
  wire [31:0] R4583;
  wire [31:0] R4582;
  wire [31:0] R4581;
  wire [31:0] R4580;
  wire [31:0] R4579;
  wire [31:0] R4578;
  wire [31:0] R4577;
  wire [31:0] R4576;
  wire [31:0] R4575;
  wire [31:0] R4574;
  wire [31:0] R4573;
  wire [31:0] R4572;
  wire [31:0] R4571;
  wire [31:0] R4570;
  wire [31:0] R4569;
  wire [31:0] R4568;
  wire [31:0] R4567;
  wire [31:0] R4566;
  wire [31:0] R4565;
  wire [31:0] R4564;
  wire [31:0] R4563;
  wire [31:0] R4562;
  wire [31:0] R4561;
  wire [31:0] R4560;
  wire [31:0] R4559;
  wire [31:0] R4558;
  wire [31:0] R4557;
  wire [31:0] R4556;
  wire [31:0] R4555;
  wire [31:0] R4554;
  wire [31:0] R4553;
  wire [31:0] R4552;
  wire [31:0] R4551;
  wire [31:0] R4550;
  wire [31:0] R4549;
  wire [31:0] R4548;
  wire [31:0] R4547;
  wire [31:0] R4546;
  wire [31:0] R4545;
  wire [31:0] R4544;
  wire [31:0] R4543;
  wire [31:0] R4542;
  wire [31:0] R4541;
  wire [31:0] R4540;
  wire [31:0] R4539;
  wire [31:0] R4538;
  wire [31:0] R4537;
  wire [31:0] R4536;
  wire [31:0] R4535;
  wire [31:0] R4534;
  wire [31:0] R4533;
  wire [31:0] R4532;
  wire [31:0] R4531;
  wire [31:0] R4530;
  wire [31:0] R4529;
  wire [31:0] R4528;
  wire [31:0] R4527;
  wire [31:0] R4526;
  wire [31:0] R4525;
  wire [31:0] R4524;
  wire [31:0] R4523;
  wire [31:0] R4522;
  wire [31:0] R4521;
  wire [31:0] R4520;
  wire [31:0] R4519;
  wire [31:0] R4518;
  wire [31:0] R4517;
  wire [31:0] R4516;
  wire [31:0] R4515;
  wire [31:0] R4514;
  wire [31:0] R4513;
  wire [31:0] R4512;
  wire [31:0] R4511;
  wire [31:0] R4510;
  wire [31:0] R4509;
  wire [31:0] R4508;
  wire [31:0] R4507;
  wire [31:0] R4506;
  wire [31:0] R4505;
  wire [31:0] R4504;
  wire [31:0] R4503;
  wire [31:0] R4502;
  wire [31:0] R4501;
  wire [31:0] R4500;
  wire [31:0] R4499;
  wire [31:0] R4498;
  wire [31:0] R4497;
  wire [31:0] R4496;
  wire [31:0] R4495;
  wire [31:0] R4494;
  wire [31:0] R4493;
  wire [31:0] R4492;
  wire [31:0] R4491;
  wire [31:0] R4490;
  wire [31:0] R4489;
  wire [31:0] R4488;
  wire [31:0] R4487;
  wire [31:0] R4486;
  wire [31:0] R4485;
  wire [31:0] R4484;
  wire [31:0] R4483;
  wire [31:0] R4482;
  wire [31:0] R4481;
  wire [31:0] R4480;
  wire [31:0] R4479;
  wire [31:0] R4478;
  wire [31:0] R4477;
  wire [31:0] R4476;
  wire [31:0] R4475;
  wire [31:0] R4474;
  wire [31:0] R4473;
  wire [31:0] R4472;
  wire [31:0] R4471;
  wire [31:0] R4470;
  wire [31:0] R4469;
  wire [31:0] R4468;
  wire [31:0] R4467;
  wire [31:0] R4466;
  wire [31:0] R4465;
  wire [31:0] R4464;
  wire [31:0] R4463;
  wire [31:0] R4462;
  wire [31:0] R4461;
  wire [31:0] R4460;
  wire [31:0] R4459;
  wire [31:0] R4458;
  wire [31:0] R4457;
  wire [31:0] R4456;
  wire [31:0] R4455;
  wire [31:0] R4454;
  wire [31:0] R4453;
  wire [31:0] R4452;
  wire [31:0] R4451;
  wire [63:0] R4450;
  wire [63:0] R4449;
  wire [63:0] R4448;
  wire [31:0] R4447;
  wire [31:0] R4446;
  wire [31:0] R4445;
  wire [31:0] R4444;
  wire [31:0] R4443;
  wire [31:0] R4442;
  wire [31:0] R4441;
  wire [31:0] R4440;
  wire [31:0] R4439;
  wire [31:0] R4438;
  wire [31:0] R4437;
  wire [31:0] R4436;
  wire [31:0] R4435;
  wire [31:0] R4434;
  wire [31:0] R4433;
  wire [31:0] R4432;
  wire [31:0] R4431;
  wire [31:0] R4430;
  wire [31:0] R4429;
  wire [31:0] R4428;
  wire [31:0] R4427;
  wire [31:0] R4426;
  wire [31:0] R4425;
  wire [31:0] R4424;
  wire [31:0] R4423;
  wire [31:0] R4422;
  wire [31:0] R4421;
  wire [31:0] R4420;
  wire [31:0] R4419;
  wire [31:0] R4418;
  wire [31:0] R4417;
  wire [31:0] R4416;
  wire [31:0] R4415;
  wire [31:0] R4414;
  wire [31:0] R4413;
  wire [31:0] R4412;
  wire [31:0] R4411;
  wire [31:0] R4410;
  wire [31:0] R4409;
  wire [31:0] R4408;
  wire [31:0] R4407;
  wire [31:0] R4406;
  wire [31:0] R4405;
  wire [31:0] R4404;
  wire [31:0] R4403;
  wire [31:0] R4402;
  wire [31:0] R4401;
  wire [31:0] R4400;
  wire [31:0] R4399;
  wire [31:0] R4398;
  wire [31:0] R4397;
  wire [31:0] R4396;
  wire [31:0] R4395;
  wire [31:0] R4394;
  wire [31:0] R4393;
  wire [31:0] R4392;
  wire [31:0] R4391;
  wire [31:0] R4390;
  wire [31:0] R4389;
  wire [31:0] R4388;
  wire [31:0] R4387;
  wire [31:0] R4386;
  wire [31:0] R4385;
  wire [31:0] R4384;
  wire [31:0] R4383;
  wire [31:0] R4382;
  wire [31:0] R4381;
  wire [31:0] R4380;
  wire [31:0] R4379;
  wire [31:0] R4378;
  wire [31:0] R4377;
  wire [31:0] R4376;
  wire [31:0] R4375;
  wire [31:0] R4374;
  wire [31:0] R4373;
  wire [31:0] R4372;
  wire [31:0] R4371;
  wire [31:0] R4370;
  wire [31:0] R4369;
  wire [31:0] R4368;
  wire [31:0] R4367;
  wire [31:0] R4366;
  wire [31:0] R4365;
  wire [31:0] R4364;
  wire [31:0] R4363;
  wire [31:0] R4362;
  wire [31:0] R4361;
  wire [31:0] R4360;
  wire [31:0] R4359;
  wire [31:0] R4358;
  wire [31:0] R4357;
  wire [31:0] R4356;
  wire [31:0] R4355;
  wire [31:0] R4354;
  wire [31:0] R4353;
  wire [31:0] R4352;
  wire [31:0] R4351;
  wire [31:0] R4350;
  wire [31:0] R4349;
  wire [31:0] R4348;
  wire [31:0] R4347;
  wire [31:0] R4346;
  wire [31:0] R4345;
  wire [31:0] R4344;
  wire [31:0] R4343;
  wire [31:0] R4342;
  wire [31:0] R4341;
  wire [31:0] R4340;
  wire [31:0] R4339;
  wire [31:0] R4338;
  wire [31:0] R4337;
  wire [31:0] R4336;
  wire [31:0] R4335;
  wire [31:0] R4334;
  wire [31:0] R4333;
  wire [31:0] R4332;
  wire [31:0] R4331;
  wire [31:0] R4330;
  wire [31:0] R4329;
  wire [31:0] R4328;
  wire [31:0] R4327;
  wire [31:0] R4326;
  wire [31:0] R4325;
  wire [31:0] R4324;
  wire [31:0] R4323;
  wire [31:0] R4322;
  wire [31:0] R4321;
  wire [31:0] R4320;
  wire [31:0] R4319;
  wire [31:0] R4318;
  wire [31:0] R4317;
  wire [31:0] R4316;
  wire [31:0] R4315;
  wire [31:0] R4314;
  wire [31:0] R4313;
  wire [31:0] R4312;
  wire [31:0] R4311;
  wire [31:0] R4310;
  wire [31:0] R4309;
  wire [31:0] R4308;
  wire [31:0] R4307;
  wire [31:0] R4306;
  wire [31:0] R4305;
  wire [31:0] R4304;
  wire [31:0] R4303;
  wire [31:0] R4302;
  wire [31:0] R4301;
  wire [31:0] R4300;
  wire [31:0] R4299;
  wire [31:0] R4298;
  wire [31:0] R4297;
  wire [31:0] R4296;
  wire [31:0] R4295;
  wire [31:0] R4294;
  wire [31:0] R4293;
  wire [31:0] R4292;
  wire [31:0] R4291;
  wire [31:0] R4290;
  wire [31:0] R4289;
  wire [31:0] R4288;
  wire [31:0] R4287;
  wire [31:0] R4286;
  wire [31:0] R4285;
  wire [31:0] R4284;
  wire [31:0] R4283;
  wire [31:0] R4282;
  wire [31:0] R4281;
  wire [31:0] R4280;
  wire [31:0] R4279;
  wire [31:0] R4278;
  wire [31:0] R4277;
  wire [31:0] R4276;
  wire [31:0] R4275;
  wire [31:0] R4274;
  wire [31:0] R4273;
  wire [31:0] R4272;
  wire [31:0] R4271;
  wire [31:0] R4270;
  wire [31:0] R4269;
  wire [31:0] R4268;
  wire [31:0] R4267;
  wire [31:0] R4266;
  wire [31:0] R4265;
  wire [31:0] R4264;
  wire [31:0] R4263;
  wire [31:0] R4262;
  wire [31:0] R4261;
  wire [31:0] R4260;
  wire [31:0] R4259;
  wire [31:0] R4258;
  wire [31:0] R4257;
  wire [31:0] R4256;
  wire [31:0] R4255;
  wire [31:0] R4254;
  wire [31:0] R4253;
  wire [31:0] R4252;
  wire [31:0] R4251;
  wire [31:0] R4250;
  wire [31:0] R4249;
  wire [31:0] R4248;
  wire [31:0] R4247;
  wire [31:0] R4246;
  wire [31:0] R4245;
  wire [31:0] R4244;
  wire [31:0] R4243;
  wire [31:0] R4242;
  wire [31:0] R4241;
  wire [31:0] R4240;
  wire [31:0] R4239;
  wire [31:0] R4238;
  wire [31:0] R4237;
  wire [31:0] R4236;
  wire [31:0] R4235;
  wire [31:0] R4234;
  wire [31:0] R4233;
  wire [31:0] R4232;
  wire [31:0] R4231;
  wire [31:0] R4230;
  wire [31:0] R4229;
  wire [31:0] R4228;
  wire [31:0] R4227;
  wire [31:0] R4226;
  wire [31:0] R4225;
  wire [31:0] R4224;
  wire [31:0] R4223;
  wire [31:0] R4222;
  wire [31:0] R4221;
  wire [31:0] R4220;
  wire [31:0] R4219;
  wire [31:0] R4218;
  wire [31:0] R4217;
  wire [31:0] R4216;
  wire [31:0] R4215;
  wire [31:0] R4214;
  wire [31:0] R4213;
  wire [31:0] R4212;
  wire [31:0] R4211;
  wire [31:0] R4210;
  wire [31:0] R4209;
  wire [31:0] R4208;
  wire [31:0] R4207;
  wire [31:0] R4206;
  wire [31:0] R4205;
  wire [31:0] R4204;
  wire [31:0] R4203;
  wire [31:0] R4202;
  wire [15:0] R4201;
  wire [63:0] R4200;
  wire [63:0] R4199;
  wire [0:0] R4198;
  wire [0:0] R4197;
  wire [0:0] R4196;
  wire [0:0] R4195;
  wire [0:0] R4194;
  wire [0:0] R4193;
  wire [0:0] R4192;
  wire [0:0] R4191;
  wire [0:0] R4190;
  wire [0:0] R4189;
  wire [0:0] R4188;
  wire [0:0] R4187;
  wire [0:0] R4186;
  wire [0:0] R4185;
  wire [0:0] R4184;
  wire [0:0] R4183;
  wire [0:0] R4182;
  wire [0:0] R4181;
  wire [0:0] R4180;
  wire [0:0] R4179;
  wire [0:0] R4178;
  wire [0:0] R4177;
  wire [0:0] R4176;
  wire [0:0] R4175;
  wire [0:0] R4174;
  wire [0:0] R4173;
  wire [0:0] R4172;
  wire [0:0] R4171;
  wire [0:0] R4170;
  wire [0:0] R4169;
  wire [0:0] R4168;
  wire [0:0] R4167;
  wire [0:0] R4166;
  wire [0:0] R4165;
  wire [0:0] R4164;
  wire [0:0] R4163;
  wire [0:0] R4162;
  wire [0:0] R4161;
  wire [0:0] R4160;
  wire [0:0] R4159;
  wire [0:0] R4158;
  wire [0:0] R4157;
  wire [0:0] R4156;
  wire [0:0] R4155;
  wire [0:0] R4154;
  wire [0:0] R4153;
  wire [0:0] R4152;
  wire [0:0] R4151;
  wire [0:0] R4150;
  wire [0:0] R4149;
  wire [0:0] R4148;
  wire [0:0] R4147;
  wire [0:0] R4146;
  wire [0:0] R4145;
  wire [0:0] R4144;
  wire [0:0] R4143;
  wire [0:0] R4142;
  wire [0:0] R4141;
  wire [0:0] R4140;
  wire [0:0] R4139;
  wire [0:0] R4138;
  wire [0:0] R4137;
  wire [0:0] R4136;
  wire [0:0] R4135;
  wire [0:0] R4134;
  wire [0:0] R4133;
  wire [0:0] R4132;
  wire [0:0] R4131;
  wire [0:0] R4130;
  wire [0:0] R4129;
  wire [0:0] R4128;
  wire [0:0] R4127;
  wire [0:0] R4126;
  wire [0:0] R4125;
  wire [0:0] R4124;
  wire [0:0] R4123;
  wire [0:0] R4122;
  wire [0:0] R4121;
  wire [0:0] R4120;
  wire [0:0] R4119;
  wire [0:0] R4118;
  wire [0:0] R4117;
  wire [0:0] R4116;
  wire [0:0] R4115;
  wire [0:0] R4114;
  wire [0:0] R4113;
  wire [0:0] R4112;
  wire [0:0] R4111;
  wire [0:0] R4110;
  wire [0:0] R4109;
  wire [0:0] R4108;
  wire [0:0] R4107;
  wire [0:0] R4106;
  wire [0:0] R4105;
  wire [0:0] R4104;
  wire [0:0] R4103;
  wire [0:0] R4102;
  wire [0:0] R4101;
  wire [0:0] R4100;
  wire [0:0] R4099;
  wire [0:0] R4098;
  wire [0:0] R4097;
  wire [0:0] R4096;
  wire [0:0] R4095;
  wire [0:0] R4094;
  wire [0:0] R4093;
  wire [0:0] R4092;
  wire [0:0] R4091;
  wire [0:0] R4090;
  wire [0:0] R4089;
  wire [0:0] R4088;
  wire [0:0] R4087;
  wire [0:0] R4086;
  wire [0:0] R4085;
  wire [0:0] R4084;
  wire [0:0] R4083;
  wire [0:0] R4082;
  wire [0:0] R4081;
  wire [0:0] R4080;
  wire [0:0] R4079;
  wire [0:0] R4078;
  wire [0:0] R4077;
  wire [0:0] R4076;
  wire [0:0] R4075;
  wire [0:0] R4074;
  wire [0:0] R4073;
  wire [0:0] R4072;
  wire [0:0] R4071;
  wire [0:0] R4070;
  wire [0:0] R4069;
  wire [0:0] R4068;
  wire [0:0] R4067;
  wire [0:0] R4066;
  wire [0:0] R4065;
  wire [0:0] R4064;
  wire [0:0] R4063;
  wire [0:0] R4062;
  wire [0:0] R4061;
  wire [0:0] R4060;
  wire [0:0] R4059;
  wire [0:0] R4058;
  wire [0:0] R4057;
  wire [0:0] R4056;
  wire [0:0] R4055;
  wire [0:0] R4054;
  wire [0:0] R4053;
  wire [0:0] R4052;
  wire [0:0] R4051;
  wire [0:0] R4050;
  wire [0:0] R4049;
  wire [0:0] R4048;
  wire [0:0] R4047;
  wire [0:0] R4046;
  wire [0:0] R4045;
  wire [0:0] R4044;
  wire [0:0] R4043;
  wire [0:0] R4042;
  wire [0:0] R4041;
  wire [0:0] R4040;
  wire [0:0] R4039;
  wire [0:0] R4038;
  wire [0:0] R4037;
  wire [0:0] R4036;
  wire [0:0] R4035;
  wire [0:0] R4034;
  wire [0:0] R4033;
  wire [0:0] R4032;
  wire [0:0] R4031;
  wire [0:0] R4030;
  wire [0:0] R4029;
  wire [0:0] R4028;
  wire [0:0] R4027;
  wire [0:0] R4026;
  wire [0:0] R4025;
  wire [0:0] R4024;
  wire [0:0] R4023;
  wire [0:0] R4022;
  wire [0:0] R4021;
  wire [0:0] R4020;
  wire [0:0] R4019;
  wire [0:0] R4018;
  wire [0:0] R4017;
  wire [0:0] R4016;
  wire [0:0] R4015;
  wire [0:0] R4014;
  wire [0:0] R4013;
  wire [0:0] R4012;
  wire [0:0] R4011;
  wire [0:0] R4010;
  wire [0:0] R4009;
  wire [0:0] R4008;
  wire [0:0] R4007;
  wire [0:0] R4006;
  wire [0:0] R4005;
  wire [0:0] R4004;
  wire [0:0] R4003;
  wire [0:0] R4002;
  wire [0:0] R4001;
  wire [0:0] R4000;
  wire [0:0] R3999;
  wire [0:0] R3998;
  wire [0:0] R3997;
  wire [0:0] R3996;
  wire [0:0] R3995;
  wire [0:0] R3994;
  wire [0:0] R3993;
  wire [0:0] R3992;
  wire [0:0] R3991;
  wire [0:0] R3990;
  wire [0:0] R3989;
  wire [0:0] R3988;
  wire [0:0] R3987;
  wire [0:0] R3986;
  wire [0:0] R3985;
  wire [0:0] R3984;
  wire [0:0] R3983;
  wire [0:0] R3982;
  wire [0:0] R3981;
  wire [0:0] R3980;
  wire [0:0] R3979;
  wire [0:0] R3978;
  wire [0:0] R3977;
  wire [0:0] R3976;
  wire [0:0] R3975;
  wire [0:0] R3974;
  wire [0:0] R3973;
  wire [0:0] R3972;
  wire [0:0] R3971;
  wire [0:0] R3970;
  wire [0:0] R3969;
  wire [0:0] R3968;
  wire [0:0] R3967;
  wire [0:0] R3966;
  wire [0:0] R3965;
  wire [0:0] R3964;
  wire [0:0] R3963;
  wire [0:0] R3962;
  wire [0:0] R3961;
  wire [0:0] R3960;
  wire [0:0] R3959;
  wire [0:0] R3958;
  wire [0:0] R3957;
  wire [0:0] R3956;
  wire [0:0] R3955;
  wire [0:0] R3954;
  wire [0:0] R3953;
  wire [0:0] R3952;
  wire [0:0] R3951;
  wire [0:0] R3950;
  wire [0:0] R3949;
  wire [0:0] R3948;
  wire [0:0] R3947;
  wire [0:0] R3946;
  wire [0:0] R3945;
  wire [0:0] R3944;
  wire [15:0] R3943;
  wire [63:0] R3942;
  wire [63:0] R3941;
  wire [31:0] R3940;
  wire [31:0] R3939;
  wire [31:0] R3938;
  wire [31:0] R3937;
  wire [31:0] R3936;
  wire [31:0] R3935;
  wire [31:0] R3934;
  wire [31:0] R3933;
  wire [31:0] R3932;
  wire [31:0] R3931;
  wire [31:0] R3930;
  wire [31:0] R3929;
  wire [31:0] R3928;
  wire [31:0] R3927;
  wire [31:0] R3926;
  wire [31:0] R3925;
  wire [31:0] R3924;
  wire [31:0] R3923;
  wire [31:0] R3922;
  wire [31:0] R3921;
  wire [31:0] R3920;
  wire [31:0] R3919;
  wire [31:0] R3918;
  wire [31:0] R3917;
  wire [31:0] R3916;
  wire [31:0] R3915;
  wire [31:0] R3914;
  wire [31:0] R3913;
  wire [31:0] R3912;
  wire [31:0] R3911;
  wire [31:0] R3910;
  wire [31:0] R3909;
  wire [31:0] R3908;
  wire [31:0] R3907;
  wire [31:0] R3906;
  wire [31:0] R3905;
  wire [31:0] R3904;
  wire [31:0] R3903;
  wire [31:0] R3902;
  wire [31:0] R3901;
  wire [31:0] R3900;
  wire [31:0] R3899;
  wire [31:0] R3898;
  wire [31:0] R3897;
  wire [31:0] R3896;
  wire [31:0] R3895;
  wire [31:0] R3894;
  wire [31:0] R3893;
  wire [31:0] R3892;
  wire [31:0] R3891;
  wire [31:0] R3890;
  wire [31:0] R3889;
  wire [31:0] R3888;
  wire [31:0] R3887;
  wire [31:0] R3886;
  wire [31:0] R3885;
  wire [31:0] R3884;
  wire [31:0] R3883;
  wire [31:0] R3882;
  wire [31:0] R3881;
  wire [31:0] R3880;
  wire [31:0] R3879;
  wire [31:0] R3878;
  wire [31:0] R3877;
  wire [31:0] R3876;
  wire [31:0] R3875;
  wire [31:0] R3874;
  wire [31:0] R3873;
  wire [31:0] R3872;
  wire [31:0] R3871;
  wire [31:0] R3870;
  wire [31:0] R3869;
  wire [31:0] R3868;
  wire [31:0] R3867;
  wire [31:0] R3866;
  wire [31:0] R3865;
  wire [31:0] R3864;
  wire [31:0] R3863;
  wire [31:0] R3862;
  wire [31:0] R3861;
  wire [31:0] R3860;
  wire [31:0] R3859;
  wire [31:0] R3858;
  wire [31:0] R3857;
  wire [31:0] R3856;
  wire [31:0] R3855;
  wire [31:0] R3854;
  wire [31:0] R3853;
  wire [31:0] R3852;
  wire [31:0] R3851;
  wire [31:0] R3850;
  wire [31:0] R3849;
  wire [31:0] R3848;
  wire [31:0] R3847;
  wire [31:0] R3846;
  wire [31:0] R3845;
  wire [31:0] R3844;
  wire [31:0] R3843;
  wire [31:0] R3842;
  wire [31:0] R3841;
  wire [31:0] R3840;
  wire [31:0] R3839;
  wire [31:0] R3838;
  wire [31:0] R3837;
  wire [31:0] R3836;
  wire [31:0] R3835;
  wire [31:0] R3834;
  wire [31:0] R3833;
  wire [31:0] R3832;
  wire [31:0] R3831;
  wire [31:0] R3830;
  wire [31:0] R3829;
  wire [31:0] R3828;
  wire [31:0] R3827;
  wire [31:0] R3826;
  wire [31:0] R3825;
  wire [31:0] R3824;
  wire [31:0] R3823;
  wire [31:0] R3822;
  wire [31:0] R3821;
  wire [31:0] R3820;
  wire [31:0] R3819;
  wire [31:0] R3818;
  wire [31:0] R3817;
  wire [31:0] R3816;
  wire [31:0] R3815;
  wire [31:0] R3814;
  wire [31:0] R3813;
  wire [31:0] R3812;
  wire [31:0] R3811;
  wire [31:0] R3810;
  wire [31:0] R3809;
  wire [31:0] R3808;
  wire [31:0] R3807;
  wire [31:0] R3806;
  wire [31:0] R3805;
  wire [31:0] R3804;
  wire [31:0] R3803;
  wire [31:0] R3802;
  wire [31:0] R3801;
  wire [31:0] R3800;
  wire [31:0] R3799;
  wire [31:0] R3798;
  wire [31:0] R3797;
  wire [31:0] R3796;
  wire [31:0] R3795;
  wire [31:0] R3794;
  wire [31:0] R3793;
  wire [31:0] R3792;
  wire [31:0] R3791;
  wire [31:0] R3790;
  wire [31:0] R3789;
  wire [31:0] R3788;
  wire [31:0] R3787;
  wire [31:0] R3786;
  wire [31:0] R3785;
  wire [31:0] R3784;
  wire [31:0] R3783;
  wire [31:0] R3782;
  wire [31:0] R3781;
  wire [31:0] R3780;
  wire [31:0] R3779;
  wire [31:0] R3778;
  wire [31:0] R3777;
  wire [31:0] R3776;
  wire [31:0] R3775;
  wire [31:0] R3774;
  wire [31:0] R3773;
  wire [31:0] R3772;
  wire [31:0] R3771;
  wire [31:0] R3770;
  wire [31:0] R3769;
  wire [31:0] R3768;
  wire [31:0] R3767;
  wire [31:0] R3766;
  wire [31:0] R3765;
  wire [31:0] R3764;
  wire [31:0] R3763;
  wire [31:0] R3762;
  wire [31:0] R3761;
  wire [31:0] R3760;
  wire [31:0] R3759;
  wire [31:0] R3758;
  wire [31:0] R3757;
  wire [31:0] R3756;
  wire [31:0] R3755;
  wire [31:0] R3754;
  wire [31:0] R3753;
  wire [31:0] R3752;
  wire [31:0] R3751;
  wire [31:0] R3750;
  wire [31:0] R3749;
  wire [31:0] R3748;
  wire [31:0] R3747;
  wire [31:0] R3746;
  wire [31:0] R3745;
  wire [31:0] R3744;
  wire [31:0] R3743;
  wire [31:0] R3742;
  wire [31:0] R3741;
  wire [31:0] R3740;
  wire [31:0] R3739;
  wire [31:0] R3738;
  wire [31:0] R3737;
  wire [31:0] R3736;
  wire [31:0] R3735;
  wire [31:0] R3734;
  wire [31:0] R3733;
  wire [31:0] R3732;
  wire [31:0] R3731;
  wire [31:0] R3730;
  wire [31:0] R3729;
  wire [31:0] R3728;
  wire [31:0] R3727;
  wire [31:0] R3726;
  wire [31:0] R3725;
  wire [31:0] R3724;
  wire [31:0] R3723;
  wire [31:0] R3722;
  wire [31:0] R3721;
  wire [31:0] R3720;
  wire [31:0] R3719;
  wire [31:0] R3718;
  wire [31:0] R3717;
  wire [31:0] R3716;
  wire [31:0] R3715;
  wire [31:0] R3714;
  wire [31:0] R3713;
  wire [31:0] R3712;
  wire [31:0] R3711;
  wire [31:0] R3710;
  wire [31:0] R3709;
  wire [31:0] R3708;
  wire [31:0] R3707;
  wire [31:0] R3706;
  wire [31:0] R3705;
  wire [31:0] R3704;
  wire [31:0] R3703;
  wire [31:0] R3702;
  wire [31:0] R3701;
  wire [31:0] R3700;
  wire [31:0] R3699;
  wire [31:0] R3698;
  wire [31:0] R3697;
  wire [31:0] R3696;
  wire [31:0] R3695;
  wire [31:0] R3694;
  wire [31:0] R3693;
  wire [31:0] R3692;
  wire [31:0] R3691;
  wire [31:0] R3690;
  wire [31:0] R3689;
  wire [31:0] R3688;
  wire [31:0] R3687;
  wire [31:0] R3686;
  wire [31:0] R3685;
  wire [31:0] R3684;
  wire [7:0] mux37;
  wire [7:0] mux36;
  wire [7:0] mux35;
  wire [7:0] mux34;
  wire [7:0] mux33;
  wire [7:0] mux32;
  wire [7:0] mux31;
  wire [7:0] mux30;
  wire [7:0] mux29;
  wire [7:0] mux28;
  wire [7:0] mux27;
  wire [7:0] mux26;
  wire [7:0] mux25;
  wire [7:0] mux24;
  wire [7:0] mux23;
  wire [7:0] mux22;
  wire [7:0] mux21;
  wire [7:0] mux20;
  wire [7:0] mux19;
  wire [7:0] mux18;
  wire [7:0] mux17;
  wire [7:0] mux16;
  wire [7:0] mux15;
  wire [7:0] mux14;
  wire [7:0] mux13;
  wire [7:0] mux12;
  wire [7:0] mux11;
  wire [7:0] mux10;
  wire [7:0] mux9;
  wire [7:0] mux8;
  wire [7:0] mux7;
  wire [7:0] mux6;
  wire [7:0] mux5;
  wire [7:0] mux4;
  wire [7:0] mux3;
  wire [7:0] mux2;
  wire [7:0] mux1;
  wire [7:0] mux0;
  wire [7:0] _3535;
  wire [63:0] _3528;
  wire [63:0] _3527;
  wire [7:0] _3688;
  wire [7:0] _3543;
  wire [63:0] _3526;
  wire [63:0] _3525;
  wire [31:0] n_idx_3541;
  wire [31:0] _3524;
  wire [31:0] _3523;
  wire [63:0] _3522;
  wire [63:0] _3521;
  wire [63:0] _3520;
  wire [63:0] _3519;
  wire [63:0] _3518;
  wire [63:0] _3517;
  wire [63:0] _3516;
  wire [63:0] _3515;
  wire [63:0] _3514;
  wire [63:0] _3513;
  wire [63:0] _3512;
  wire [63:0] _3511;
  wire [63:0] _3510;
  wire [63:0] _3509;
  wire [63:0] _3508;
  wire [63:0] _3507;
  wire [63:0] _3506;
  wire [63:0] _3505;
  wire [63:0] _3504;
  wire [63:0] _3503;
  wire [63:0] _3502;
  wire [63:0] _3501;
  wire [63:0] _3500;
  wire [63:0] _3499;
  wire [63:0] _3498;
  wire [63:0] _3497;
  wire [63:0] _3496;
  wire [63:0] _3495;
  wire [63:0] _3494;
  wire [63:0] _3493;
  wire [63:0] _3492;
  wire [63:0] _3491;
  wire [63:0] _3490;
  wire [63:0] _3489;
  wire [63:0] _3488;
  wire [63:0] _3487;
  wire [63:0] _3486;
  wire [63:0] _3485;
  wire [63:0] _3484;
  wire [63:0] _3483;
  wire [63:0] _3482;
  wire [63:0] _3481;
  wire [63:0] _3480;
  wire [63:0] _3479;
  wire [63:0] _3478;
  wire [63:0] _3477;
  wire [63:0] _3476;
  wire [63:0] _3475;
  wire [63:0] _3474;
  wire [63:0] _3473;
  wire [63:0] _3472;
  wire [63:0] _3471;
  wire [63:0] _3470;
  wire [63:0] _3469;
  wire [63:0] _3468;
  wire [63:0] _3467;
  wire [63:0] _3466;
  wire [63:0] _3465;
  wire [63:0] _3464;
  wire [63:0] _3463;
  wire [63:0] _3462;
  wire [63:0] _3461;
  wire [63:0] _3460;
  wire [63:0] _3459;
  wire [63:0] _3458;
  wire [63:0] _3457;
  wire [63:0] _3456;
  wire [63:0] _3455;
  wire [63:0] _3454;
  wire [63:0] _3453;
  wire [63:0] _3452;
  wire [63:0] _3451;
  wire [63:0] _3450;
  wire [63:0] _3449;
  wire [63:0] _3448;
  wire [63:0] _3447;
  wire [63:0] _3446;
  wire [63:0] _3445;
  wire [63:0] _3444;
  wire [63:0] _3443;
  wire [63:0] _3442;
  wire [31:0] _3441;
  wire [63:0] _3440;
  wire [63:0] _3439;
  wire [63:0] _3438;
  wire [0:0] ifout3549;
  wire [63:0] _3437;
  wire [63:0] _3436;
  wire [63:0] _3435;
  wire [63:0] _3434;
  wire [63:0] _3433;
  wire [63:0] _3432;
  wire [7:0] _3551;
  wire [63:0] _3431;
  wire [63:0] _3430;
  wire [31:0] n_idx_3550;
  wire [31:0] _3429;
  wire [31:0] _3428;
  wire [63:0] _3427;
  wire [63:0] _3426;
  wire [63:0] _3425;
  wire [63:0] _3424;
  wire [63:0] _3423;
  wire [63:0] _3422;
  wire [63:0] _3421;
  wire [63:0] _3420;
  wire [63:0] _3419;
  wire [63:0] _3418;
  wire [63:0] _3417;
  wire [63:0] _3416;
  wire [63:0] _3415;
  wire [63:0] _3414;
  wire [63:0] _3413;
  wire [63:0] _3412;
  wire [63:0] _3411;
  wire [63:0] _3410;
  wire [63:0] _3409;
  wire [63:0] _3408;
  wire [63:0] _3407;
  wire [63:0] _3406;
  wire [63:0] _3405;
  wire [63:0] _3404;
  wire [63:0] _3403;
  wire [63:0] _3402;
  wire [63:0] _3401;
  wire [63:0] _3400;
  wire [63:0] _3399;
  wire [63:0] _3398;
  wire [63:0] _3397;
  wire [63:0] _3396;
  wire [63:0] _3395;
  wire [63:0] _3394;
  wire [63:0] _3393;
  wire [63:0] _3392;
  wire [63:0] _3391;
  wire [63:0] _3390;
  wire [63:0] _3389;
  wire [63:0] _3388;
  wire [63:0] _3387;
  wire [63:0] _3386;
  wire [63:0] _3385;
  wire [63:0] _3384;
  wire [63:0] _3383;
  wire [63:0] _3382;
  wire [63:0] _3381;
  wire [63:0] _3380;
  wire [63:0] _3379;
  wire [63:0] _3378;
  wire [63:0] _3377;
  wire [63:0] _3376;
  wire [63:0] _3375;
  wire [63:0] _3374;
  wire [63:0] _3373;
  wire [63:0] _3372;
  wire [63:0] _3371;
  wire [63:0] _3370;
  wire [63:0] _3369;
  wire [63:0] _3368;
  wire [63:0] _3367;
  wire [63:0] _3366;
  wire [63:0] _3365;
  wire [63:0] _3364;
  wire [63:0] _3363;
  wire [63:0] _3362;
  wire [63:0] _3361;
  wire [63:0] _3360;
  wire [63:0] _3359;
  wire [63:0] _3358;
  wire [63:0] _3357;
  wire [63:0] _3356;
  wire [63:0] _3355;
  wire [63:0] _3354;
  wire [63:0] _3353;
  wire [63:0] _3352;
  wire [63:0] _3351;
  wire [63:0] _3350;
  wire [63:0] _3349;
  wire [63:0] _3348;
  wire [63:0] _3347;
  wire [31:0] _3346;
  wire [63:0] _3345;
  wire [63:0] _3344;
  wire [63:0] _3343;
  wire [0:0] ifout3451;
  wire [63:0] _3342;
  wire [63:0] _3341;
  wire [63:0] _3340;
  wire [63:0] _3339;
  wire [63:0] _3338;
  wire [63:0] _3337;
  wire [7:0] _3559;
  wire [63:0] _3336;
  wire [63:0] _3335;
  wire [31:0] n_idx_3558;
  wire [31:0] _3334;
  wire [31:0] _3333;
  wire [63:0] _3332;
  wire [63:0] _3331;
  wire [63:0] _3330;
  wire [63:0] _3329;
  wire [63:0] _3328;
  wire [63:0] _3327;
  wire [63:0] _3326;
  wire [63:0] _3325;
  wire [63:0] _3324;
  wire [63:0] _3323;
  wire [63:0] _3322;
  wire [63:0] _3321;
  wire [63:0] _3320;
  wire [63:0] _3319;
  wire [63:0] _3318;
  wire [63:0] _3317;
  wire [63:0] _3316;
  wire [63:0] _3315;
  wire [63:0] _3314;
  wire [63:0] _3313;
  wire [63:0] _3312;
  wire [63:0] _3311;
  wire [63:0] _3310;
  wire [63:0] _3309;
  wire [63:0] _3308;
  wire [63:0] _3307;
  wire [63:0] _3306;
  wire [63:0] _3305;
  wire [63:0] _3304;
  wire [63:0] _3303;
  wire [63:0] _3302;
  wire [63:0] _3301;
  wire [63:0] _3300;
  wire [63:0] _3299;
  wire [63:0] _3298;
  wire [63:0] _3297;
  wire [63:0] _3296;
  wire [63:0] _3295;
  wire [63:0] _3294;
  wire [63:0] _3293;
  wire [63:0] _3292;
  wire [63:0] _3291;
  wire [63:0] _3290;
  wire [63:0] _3289;
  wire [63:0] _3288;
  wire [63:0] _3287;
  wire [63:0] _3286;
  wire [63:0] _3285;
  wire [63:0] _3284;
  wire [63:0] _3283;
  wire [63:0] _3282;
  wire [63:0] _3281;
  wire [63:0] _3280;
  wire [63:0] _3279;
  wire [63:0] _3278;
  wire [63:0] _3277;
  wire [63:0] _3276;
  wire [63:0] _3275;
  wire [63:0] _3274;
  wire [63:0] _3273;
  wire [63:0] _3272;
  wire [63:0] _3271;
  wire [63:0] _3270;
  wire [63:0] _3269;
  wire [63:0] _3268;
  wire [63:0] _3267;
  wire [63:0] _3266;
  wire [63:0] _3265;
  wire [63:0] _3264;
  wire [63:0] _3263;
  wire [63:0] _3262;
  wire [63:0] _3261;
  wire [63:0] _3260;
  wire [63:0] _3259;
  wire [63:0] _3258;
  wire [63:0] _3257;
  wire [63:0] _3256;
  wire [63:0] _3255;
  wire [63:0] _3254;
  wire [63:0] _3253;
  wire [63:0] _3252;
  wire [31:0] _3251;
  wire [63:0] _3250;
  wire [63:0] _3249;
  wire [63:0] _3248;
  wire [0:0] ifout3353;
  wire [63:0] _3247;
  wire [63:0] _3246;
  wire [63:0] _3245;
  wire [63:0] _3244;
  wire [63:0] _3243;
  wire [63:0] _3242;
  wire [7:0] _3567;
  wire [63:0] _3241;
  wire [63:0] _3240;
  wire [31:0] n_idx_3566;
  wire [31:0] _3239;
  wire [31:0] _3238;
  wire [63:0] _3237;
  wire [63:0] _3236;
  wire [63:0] _3235;
  wire [63:0] _3234;
  wire [63:0] _3233;
  wire [63:0] _3232;
  wire [63:0] _3231;
  wire [63:0] _3230;
  wire [63:0] _3229;
  wire [63:0] _3228;
  wire [63:0] _3227;
  wire [63:0] _3226;
  wire [63:0] _3225;
  wire [63:0] _3224;
  wire [63:0] _3223;
  wire [63:0] _3222;
  wire [63:0] _3221;
  wire [63:0] _3220;
  wire [63:0] _3219;
  wire [63:0] _3218;
  wire [63:0] _3217;
  wire [63:0] _3216;
  wire [63:0] _3215;
  wire [63:0] _3214;
  wire [63:0] _3213;
  wire [63:0] _3212;
  wire [63:0] _3211;
  wire [63:0] _3210;
  wire [63:0] _3209;
  wire [63:0] _3208;
  wire [63:0] _3207;
  wire [63:0] _3206;
  wire [63:0] _3205;
  wire [63:0] _3204;
  wire [63:0] _3203;
  wire [63:0] _3202;
  wire [63:0] _3201;
  wire [63:0] _3200;
  wire [63:0] _3199;
  wire [63:0] _3198;
  wire [63:0] _3197;
  wire [63:0] _3196;
  wire [63:0] _3195;
  wire [63:0] _3194;
  wire [63:0] _3193;
  wire [63:0] _3192;
  wire [63:0] _3191;
  wire [63:0] _3190;
  wire [63:0] _3189;
  wire [63:0] _3188;
  wire [63:0] _3187;
  wire [63:0] _3186;
  wire [63:0] _3185;
  wire [63:0] _3184;
  wire [63:0] _3183;
  wire [63:0] _3182;
  wire [63:0] _3181;
  wire [63:0] _3180;
  wire [63:0] _3179;
  wire [63:0] _3178;
  wire [63:0] _3177;
  wire [63:0] _3176;
  wire [63:0] _3175;
  wire [63:0] _3174;
  wire [63:0] _3173;
  wire [63:0] _3172;
  wire [63:0] _3171;
  wire [63:0] _3170;
  wire [63:0] _3169;
  wire [63:0] _3168;
  wire [63:0] _3167;
  wire [63:0] _3166;
  wire [63:0] _3165;
  wire [63:0] _3164;
  wire [63:0] _3163;
  wire [63:0] _3162;
  wire [63:0] _3161;
  wire [63:0] _3160;
  wire [63:0] _3159;
  wire [63:0] _3158;
  wire [63:0] _3157;
  wire [31:0] _3156;
  wire [63:0] _3155;
  wire [63:0] _3154;
  wire [63:0] _3153;
  wire [0:0] ifout3255;
  wire [63:0] _3152;
  wire [63:0] _3151;
  wire [63:0] _3150;
  wire [63:0] _3149;
  wire [63:0] _3148;
  wire [63:0] _3147;
  wire [7:0] _3575;
  wire [63:0] _3146;
  wire [63:0] _3145;
  wire [31:0] n_idx_3574;
  wire [31:0] _3144;
  wire [31:0] _3143;
  wire [63:0] _3142;
  wire [63:0] _3141;
  wire [63:0] _3140;
  wire [63:0] _3139;
  wire [63:0] _3138;
  wire [63:0] _3137;
  wire [63:0] _3136;
  wire [63:0] _3135;
  wire [63:0] _3134;
  wire [63:0] _3133;
  wire [63:0] _3132;
  wire [63:0] _3131;
  wire [63:0] _3130;
  wire [63:0] _3129;
  wire [63:0] _3128;
  wire [63:0] _3127;
  wire [63:0] _3126;
  wire [63:0] _3125;
  wire [63:0] _3124;
  wire [63:0] _3123;
  wire [63:0] _3122;
  wire [63:0] _3121;
  wire [63:0] _3120;
  wire [63:0] _3119;
  wire [63:0] _3118;
  wire [63:0] _3117;
  wire [63:0] _3116;
  wire [63:0] _3115;
  wire [63:0] _3114;
  wire [63:0] _3113;
  wire [63:0] _3112;
  wire [63:0] _3111;
  wire [63:0] _3110;
  wire [63:0] _3109;
  wire [63:0] _3108;
  wire [63:0] _3107;
  wire [63:0] _3106;
  wire [63:0] _3105;
  wire [63:0] _3104;
  wire [63:0] _3103;
  wire [63:0] _3102;
  wire [63:0] _3101;
  wire [63:0] _3100;
  wire [63:0] _3099;
  wire [63:0] _3098;
  wire [63:0] _3097;
  wire [63:0] _3096;
  wire [63:0] _3095;
  wire [63:0] _3094;
  wire [63:0] _3093;
  wire [63:0] _3092;
  wire [63:0] _3091;
  wire [63:0] _3090;
  wire [63:0] _3089;
  wire [63:0] _3088;
  wire [63:0] _3087;
  wire [63:0] _3086;
  wire [63:0] _3085;
  wire [63:0] _3084;
  wire [63:0] _3083;
  wire [63:0] _3082;
  wire [63:0] _3081;
  wire [63:0] _3080;
  wire [63:0] _3079;
  wire [63:0] _3078;
  wire [63:0] _3077;
  wire [63:0] _3076;
  wire [63:0] _3075;
  wire [63:0] _3074;
  wire [63:0] _3073;
  wire [63:0] _3072;
  wire [63:0] _3071;
  wire [63:0] _3070;
  wire [63:0] _3069;
  wire [63:0] _3068;
  wire [63:0] _3067;
  wire [63:0] _3066;
  wire [63:0] _3065;
  wire [63:0] _3064;
  wire [63:0] _3063;
  wire [63:0] _3062;
  wire [31:0] _3061;
  wire [63:0] _3060;
  wire [63:0] _3059;
  wire [63:0] _3058;
  wire [0:0] ifout3157;
  wire [63:0] _3057;
  wire [63:0] _3056;
  wire [63:0] _3055;
  wire [63:0] _3054;
  wire [63:0] _3053;
  wire [63:0] _3052;
  wire [7:0] _3583;
  wire [63:0] _3051;
  wire [63:0] _3050;
  wire [31:0] n_idx_3582;
  wire [31:0] _3049;
  wire [31:0] _3048;
  wire [63:0] _3047;
  wire [63:0] _3046;
  wire [63:0] _3045;
  wire [63:0] _3044;
  wire [63:0] _3043;
  wire [63:0] _3042;
  wire [63:0] _3041;
  wire [63:0] _3040;
  wire [63:0] _3039;
  wire [63:0] _3038;
  wire [63:0] _3037;
  wire [63:0] _3036;
  wire [63:0] _3035;
  wire [63:0] _3034;
  wire [63:0] _3033;
  wire [63:0] _3032;
  wire [63:0] _3031;
  wire [63:0] _3030;
  wire [63:0] _3029;
  wire [63:0] _3028;
  wire [63:0] _3027;
  wire [63:0] _3026;
  wire [63:0] _3025;
  wire [63:0] _3024;
  wire [63:0] _3023;
  wire [63:0] _3022;
  wire [63:0] _3021;
  wire [63:0] _3020;
  wire [63:0] _3019;
  wire [63:0] _3018;
  wire [63:0] _3017;
  wire [63:0] _3016;
  wire [63:0] _3015;
  wire [63:0] _3014;
  wire [63:0] _3013;
  wire [63:0] _3012;
  wire [63:0] _3011;
  wire [63:0] _3010;
  wire [63:0] _3009;
  wire [63:0] _3008;
  wire [63:0] _3007;
  wire [63:0] _3006;
  wire [63:0] _3005;
  wire [63:0] _3004;
  wire [63:0] _3003;
  wire [63:0] _3002;
  wire [63:0] _3001;
  wire [63:0] _3000;
  wire [63:0] _2999;
  wire [63:0] _2998;
  wire [63:0] _2997;
  wire [63:0] _2996;
  wire [63:0] _2995;
  wire [63:0] _2994;
  wire [63:0] _2993;
  wire [63:0] _2992;
  wire [63:0] _2991;
  wire [63:0] _2990;
  wire [63:0] _2989;
  wire [63:0] _2988;
  wire [63:0] _2987;
  wire [63:0] _2986;
  wire [63:0] _2985;
  wire [63:0] _2984;
  wire [63:0] _2983;
  wire [63:0] _2982;
  wire [63:0] _2981;
  wire [63:0] _2980;
  wire [63:0] _2979;
  wire [63:0] _2978;
  wire [63:0] _2977;
  wire [63:0] _2976;
  wire [63:0] _2975;
  wire [63:0] _2974;
  wire [63:0] _2973;
  wire [63:0] _2972;
  wire [63:0] _2971;
  wire [63:0] _2970;
  wire [63:0] _2969;
  wire [63:0] _2968;
  wire [63:0] _2967;
  wire [31:0] _2966;
  wire [63:0] _2965;
  wire [63:0] _2964;
  wire [63:0] _2963;
  wire [0:0] ifout3059;
  wire [63:0] _2962;
  wire [63:0] _2961;
  wire [63:0] _2960;
  wire [63:0] _2959;
  wire [63:0] _2958;
  wire [63:0] _2957;
  wire [7:0] _3591;
  wire [63:0] _2956;
  wire [63:0] _2955;
  wire [31:0] n_idx_3590;
  wire [31:0] _2954;
  wire [31:0] _2953;
  wire [63:0] _2952;
  wire [63:0] _2951;
  wire [63:0] _2950;
  wire [63:0] _2949;
  wire [63:0] _2948;
  wire [63:0] _2947;
  wire [63:0] _2946;
  wire [63:0] _2945;
  wire [63:0] _2944;
  wire [63:0] _2943;
  wire [63:0] _2942;
  wire [63:0] _2941;
  wire [63:0] _2940;
  wire [63:0] _2939;
  wire [63:0] _2938;
  wire [63:0] _2937;
  wire [63:0] _2936;
  wire [63:0] _2935;
  wire [63:0] _2934;
  wire [63:0] _2933;
  wire [63:0] _2932;
  wire [63:0] _2931;
  wire [63:0] _2930;
  wire [63:0] _2929;
  wire [63:0] _2928;
  wire [63:0] _2927;
  wire [63:0] _2926;
  wire [63:0] _2925;
  wire [63:0] _2924;
  wire [63:0] _2923;
  wire [63:0] _2922;
  wire [63:0] _2921;
  wire [63:0] _2920;
  wire [63:0] _2919;
  wire [63:0] _2918;
  wire [63:0] _2917;
  wire [63:0] _2916;
  wire [63:0] _2915;
  wire [63:0] _2914;
  wire [63:0] _2913;
  wire [63:0] _2912;
  wire [63:0] _2911;
  wire [63:0] _2910;
  wire [63:0] _2909;
  wire [63:0] _2908;
  wire [63:0] _2907;
  wire [63:0] _2906;
  wire [63:0] _2905;
  wire [63:0] _2904;
  wire [63:0] _2903;
  wire [63:0] _2902;
  wire [63:0] _2901;
  wire [63:0] _2900;
  wire [63:0] _2899;
  wire [63:0] _2898;
  wire [63:0] _2897;
  wire [63:0] _2896;
  wire [63:0] _2895;
  wire [63:0] _2894;
  wire [63:0] _2893;
  wire [63:0] _2892;
  wire [63:0] _2891;
  wire [63:0] _2890;
  wire [63:0] _2889;
  wire [63:0] _2888;
  wire [63:0] _2887;
  wire [63:0] _2886;
  wire [63:0] _2885;
  wire [63:0] _2884;
  wire [63:0] _2883;
  wire [63:0] _2882;
  wire [63:0] _2881;
  wire [63:0] _2880;
  wire [63:0] _2879;
  wire [63:0] _2878;
  wire [63:0] _2877;
  wire [63:0] _2876;
  wire [63:0] _2875;
  wire [63:0] _2874;
  wire [63:0] _2873;
  wire [63:0] _2872;
  wire [31:0] _2871;
  wire [63:0] _2870;
  wire [63:0] _2869;
  wire [63:0] _2868;
  wire [0:0] ifout2961;
  wire [63:0] _2867;
  wire [63:0] _2866;
  wire [63:0] _2865;
  wire [63:0] _2864;
  wire [63:0] _2863;
  wire [63:0] _2862;
  wire [7:0] _3599;
  wire [63:0] _2861;
  wire [63:0] _2860;
  wire [31:0] n_idx_3598;
  wire [31:0] _2859;
  wire [31:0] _2858;
  wire [63:0] _2857;
  wire [63:0] _2856;
  wire [63:0] _2855;
  wire [63:0] _2854;
  wire [63:0] _2853;
  wire [63:0] _2852;
  wire [63:0] _2851;
  wire [63:0] _2850;
  wire [63:0] _2849;
  wire [63:0] _2848;
  wire [63:0] _2847;
  wire [63:0] _2846;
  wire [63:0] _2845;
  wire [63:0] _2844;
  wire [63:0] _2843;
  wire [63:0] _2842;
  wire [63:0] _2841;
  wire [63:0] _2840;
  wire [63:0] _2839;
  wire [63:0] _2838;
  wire [63:0] _2837;
  wire [63:0] _2836;
  wire [63:0] _2835;
  wire [63:0] _2834;
  wire [63:0] _2833;
  wire [63:0] _2832;
  wire [63:0] _2831;
  wire [63:0] _2830;
  wire [63:0] _2829;
  wire [63:0] _2828;
  wire [63:0] _2827;
  wire [63:0] _2826;
  wire [63:0] _2825;
  wire [63:0] _2824;
  wire [63:0] _2823;
  wire [63:0] _2822;
  wire [63:0] _2821;
  wire [63:0] _2820;
  wire [63:0] _2819;
  wire [63:0] _2818;
  wire [63:0] _2817;
  wire [63:0] _2816;
  wire [63:0] _2815;
  wire [63:0] _2814;
  wire [63:0] _2813;
  wire [63:0] _2812;
  wire [63:0] _2811;
  wire [63:0] _2810;
  wire [63:0] _2809;
  wire [63:0] _2808;
  wire [63:0] _2807;
  wire [63:0] _2806;
  wire [63:0] _2805;
  wire [63:0] _2804;
  wire [63:0] _2803;
  wire [63:0] _2802;
  wire [63:0] _2801;
  wire [63:0] _2800;
  wire [63:0] _2799;
  wire [63:0] _2798;
  wire [63:0] _2797;
  wire [63:0] _2796;
  wire [63:0] _2795;
  wire [63:0] _2794;
  wire [63:0] _2793;
  wire [63:0] _2792;
  wire [63:0] _2791;
  wire [63:0] _2790;
  wire [63:0] _2789;
  wire [63:0] _2788;
  wire [63:0] _2787;
  wire [63:0] _2786;
  wire [63:0] _2785;
  wire [63:0] _2784;
  wire [63:0] _2783;
  wire [63:0] _2782;
  wire [63:0] _2781;
  wire [63:0] _2780;
  wire [63:0] _2779;
  wire [63:0] _2778;
  wire [63:0] _2777;
  wire [31:0] _2776;
  wire [63:0] _2775;
  wire [63:0] _2774;
  wire [63:0] _2773;
  wire [0:0] ifout2863;
  wire [63:0] _2772;
  wire [63:0] _2771;
  wire [63:0] _2770;
  wire [63:0] _2769;
  wire [63:0] _2768;
  wire [63:0] _2767;
  wire [7:0] _3608;
  wire [63:0] _2766;
  wire [63:0] _2765;
  wire [31:0] n_idx_3607;
  wire [31:0] _2764;
  wire [31:0] _2763;
  wire [63:0] _2762;
  wire [63:0] _2761;
  wire [63:0] _2760;
  wire [63:0] _2759;
  wire [63:0] _2758;
  wire [63:0] _2757;
  wire [63:0] _2756;
  wire [63:0] _2755;
  wire [63:0] _2754;
  wire [63:0] _2753;
  wire [63:0] _2752;
  wire [63:0] _2751;
  wire [63:0] _2750;
  wire [63:0] _2749;
  wire [63:0] _2748;
  wire [63:0] _2747;
  wire [63:0] _2746;
  wire [63:0] _2745;
  wire [63:0] _2744;
  wire [63:0] _2743;
  wire [63:0] _2742;
  wire [63:0] _2741;
  wire [63:0] _2740;
  wire [63:0] _2739;
  wire [63:0] _2738;
  wire [63:0] _2737;
  wire [63:0] _2736;
  wire [63:0] _2735;
  wire [63:0] _2734;
  wire [63:0] _2733;
  wire [63:0] _2732;
  wire [63:0] _2731;
  wire [63:0] _2730;
  wire [63:0] _2729;
  wire [63:0] _2728;
  wire [63:0] _2727;
  wire [63:0] _2726;
  wire [63:0] _2725;
  wire [63:0] _2724;
  wire [63:0] _2723;
  wire [63:0] _2722;
  wire [63:0] _2721;
  wire [63:0] _2720;
  wire [63:0] _2719;
  wire [63:0] _2718;
  wire [63:0] _2717;
  wire [63:0] _2716;
  wire [63:0] _2715;
  wire [63:0] _2714;
  wire [63:0] _2713;
  wire [63:0] _2712;
  wire [63:0] _2711;
  wire [63:0] _2710;
  wire [63:0] _2709;
  wire [63:0] _2708;
  wire [63:0] _2707;
  wire [63:0] _2706;
  wire [63:0] _2705;
  wire [63:0] _2704;
  wire [63:0] _2703;
  wire [63:0] _2702;
  wire [63:0] _2701;
  wire [63:0] _2700;
  wire [63:0] _2699;
  wire [63:0] _2698;
  wire [63:0] _2697;
  wire [63:0] _2696;
  wire [63:0] _2695;
  wire [63:0] _2694;
  wire [63:0] _2693;
  wire [63:0] _2692;
  wire [63:0] _2691;
  wire [63:0] _2690;
  wire [63:0] _2689;
  wire [63:0] _2688;
  wire [63:0] _2687;
  wire [63:0] _2686;
  wire [63:0] _2685;
  wire [63:0] _2684;
  wire [63:0] _2683;
  wire [63:0] _2682;
  wire [31:0] _2681;
  wire [63:0] _2680;
  wire [63:0] _2679;
  wire [63:0] _2678;
  wire [0:0] ifout2765;
  wire [63:0] _2677;
  wire [63:0] _2676;
  wire [63:0] _2675;
  wire [63:0] _2674;
  wire [63:0] _2673;
  wire [63:0] _2672;
  wire [7:0] _3616;
  wire [63:0] _2671;
  wire [63:0] _2670;
  wire [31:0] n_idx_3615;
  wire [31:0] _2669;
  wire [31:0] _2668;
  wire [63:0] _2667;
  wire [63:0] _2666;
  wire [63:0] _2665;
  wire [63:0] _2664;
  wire [63:0] _2663;
  wire [63:0] _2662;
  wire [63:0] _2661;
  wire [63:0] _2660;
  wire [63:0] _2659;
  wire [63:0] _2658;
  wire [63:0] _2657;
  wire [63:0] _2656;
  wire [63:0] _2655;
  wire [63:0] _2654;
  wire [63:0] _2653;
  wire [63:0] _2652;
  wire [63:0] _2651;
  wire [63:0] _2650;
  wire [63:0] _2649;
  wire [63:0] _2648;
  wire [63:0] _2647;
  wire [63:0] _2646;
  wire [63:0] _2645;
  wire [63:0] _2644;
  wire [63:0] _2643;
  wire [63:0] _2642;
  wire [63:0] _2641;
  wire [63:0] _2640;
  wire [63:0] _2639;
  wire [63:0] _2638;
  wire [63:0] _2637;
  wire [63:0] _2636;
  wire [63:0] _2635;
  wire [63:0] _2634;
  wire [63:0] _2633;
  wire [63:0] _2632;
  wire [63:0] _2631;
  wire [63:0] _2630;
  wire [63:0] _2629;
  wire [63:0] _2628;
  wire [63:0] _2627;
  wire [63:0] _2626;
  wire [63:0] _2625;
  wire [63:0] _2624;
  wire [63:0] _2623;
  wire [63:0] _2622;
  wire [63:0] _2621;
  wire [63:0] _2620;
  wire [63:0] _2619;
  wire [63:0] _2618;
  wire [63:0] _2617;
  wire [63:0] _2616;
  wire [63:0] _2615;
  wire [63:0] _2614;
  wire [63:0] _2613;
  wire [63:0] _2612;
  wire [63:0] _2611;
  wire [63:0] _2610;
  wire [63:0] _2609;
  wire [63:0] _2608;
  wire [63:0] _2607;
  wire [63:0] _2606;
  wire [63:0] _2605;
  wire [63:0] _2604;
  wire [63:0] _2603;
  wire [63:0] _2602;
  wire [63:0] _2601;
  wire [63:0] _2600;
  wire [63:0] _2599;
  wire [63:0] _2598;
  wire [63:0] _2597;
  wire [63:0] _2596;
  wire [63:0] _2595;
  wire [63:0] _2594;
  wire [63:0] _2593;
  wire [63:0] _2592;
  wire [63:0] _2591;
  wire [63:0] _2590;
  wire [63:0] _2589;
  wire [63:0] _2588;
  wire [63:0] _2587;
  wire [31:0] _2586;
  wire [63:0] _2585;
  wire [63:0] _2584;
  wire [63:0] _2583;
  wire [0:0] ifout2667;
  wire [63:0] _2582;
  wire [63:0] _2581;
  wire [63:0] _2580;
  wire [63:0] _2579;
  wire [63:0] _2578;
  wire [63:0] _2577;
  wire [7:0] _3624;
  wire [63:0] _2576;
  wire [63:0] _2575;
  wire [31:0] n_idx_3623;
  wire [31:0] _2574;
  wire [31:0] _2573;
  wire [63:0] _2572;
  wire [63:0] _2571;
  wire [63:0] _2570;
  wire [63:0] _2569;
  wire [63:0] _2568;
  wire [63:0] _2567;
  wire [63:0] _2566;
  wire [63:0] _2565;
  wire [63:0] _2564;
  wire [63:0] _2563;
  wire [63:0] _2562;
  wire [63:0] _2561;
  wire [63:0] _2560;
  wire [63:0] _2559;
  wire [63:0] _2558;
  wire [63:0] _2557;
  wire [63:0] _2556;
  wire [63:0] _2555;
  wire [63:0] _2554;
  wire [63:0] _2553;
  wire [63:0] _2552;
  wire [63:0] _2551;
  wire [63:0] _2550;
  wire [63:0] _2549;
  wire [63:0] _2548;
  wire [63:0] _2547;
  wire [63:0] _2546;
  wire [63:0] _2545;
  wire [63:0] _2544;
  wire [63:0] _2543;
  wire [63:0] _2542;
  wire [63:0] _2541;
  wire [63:0] _2540;
  wire [63:0] _2539;
  wire [63:0] _2538;
  wire [63:0] _2537;
  wire [63:0] _2536;
  wire [63:0] _2535;
  wire [63:0] _2534;
  wire [63:0] _2533;
  wire [63:0] _2532;
  wire [63:0] _2531;
  wire [63:0] _2530;
  wire [63:0] _2529;
  wire [63:0] _2528;
  wire [63:0] _2527;
  wire [63:0] _2526;
  wire [63:0] _2525;
  wire [63:0] _2524;
  wire [63:0] _2523;
  wire [63:0] _2522;
  wire [63:0] _2521;
  wire [63:0] _2520;
  wire [63:0] _2519;
  wire [63:0] _2518;
  wire [63:0] _2517;
  wire [63:0] _2516;
  wire [63:0] _2515;
  wire [63:0] _2514;
  wire [63:0] _2513;
  wire [63:0] _2512;
  wire [63:0] _2511;
  wire [63:0] _2510;
  wire [63:0] _2509;
  wire [63:0] _2508;
  wire [63:0] _2507;
  wire [63:0] _2506;
  wire [63:0] _2505;
  wire [63:0] _2504;
  wire [63:0] _2503;
  wire [63:0] _2502;
  wire [63:0] _2501;
  wire [63:0] _2500;
  wire [63:0] _2499;
  wire [63:0] _2498;
  wire [63:0] _2497;
  wire [63:0] _2496;
  wire [63:0] _2495;
  wire [63:0] _2494;
  wire [63:0] _2493;
  wire [63:0] _2492;
  wire [31:0] _2491;
  wire [63:0] _2490;
  wire [63:0] _2489;
  wire [63:0] _2488;
  wire [0:0] ifout2569;
  wire [63:0] _2487;
  wire [63:0] _2486;
  wire [63:0] _2485;
  wire [63:0] _2484;
  wire [63:0] _2483;
  wire [63:0] _2482;
  wire [7:0] _3632;
  wire [63:0] _2481;
  wire [63:0] _2480;
  wire [31:0] n_idx_3631;
  wire [31:0] _2479;
  wire [31:0] _2478;
  wire [63:0] _2477;
  wire [63:0] _2476;
  wire [63:0] _2475;
  wire [63:0] _2474;
  wire [63:0] _2473;
  wire [63:0] _2472;
  wire [63:0] _2471;
  wire [63:0] _2470;
  wire [63:0] _2469;
  wire [63:0] _2468;
  wire [63:0] _2467;
  wire [63:0] _2466;
  wire [63:0] _2465;
  wire [63:0] _2464;
  wire [63:0] _2463;
  wire [63:0] _2462;
  wire [63:0] _2461;
  wire [63:0] _2460;
  wire [63:0] _2459;
  wire [63:0] _2458;
  wire [63:0] _2457;
  wire [63:0] _2456;
  wire [63:0] _2455;
  wire [63:0] _2454;
  wire [63:0] _2453;
  wire [63:0] _2452;
  wire [63:0] _2451;
  wire [63:0] _2450;
  wire [63:0] _2449;
  wire [63:0] _2448;
  wire [63:0] _2447;
  wire [63:0] _2446;
  wire [63:0] _2445;
  wire [63:0] _2444;
  wire [63:0] _2443;
  wire [63:0] _2442;
  wire [63:0] _2441;
  wire [63:0] _2440;
  wire [63:0] _2439;
  wire [63:0] _2438;
  wire [63:0] _2437;
  wire [63:0] _2436;
  wire [63:0] _2435;
  wire [63:0] _2434;
  wire [63:0] _2433;
  wire [63:0] _2432;
  wire [63:0] _2431;
  wire [63:0] _2430;
  wire [63:0] _2429;
  wire [63:0] _2428;
  wire [63:0] _2427;
  wire [63:0] _2426;
  wire [63:0] _2425;
  wire [63:0] _2424;
  wire [63:0] _2423;
  wire [63:0] _2422;
  wire [63:0] _2421;
  wire [63:0] _2420;
  wire [63:0] _2419;
  wire [63:0] _2418;
  wire [63:0] _2417;
  wire [63:0] _2416;
  wire [63:0] _2415;
  wire [63:0] _2414;
  wire [63:0] _2413;
  wire [63:0] _2412;
  wire [63:0] _2411;
  wire [63:0] _2410;
  wire [63:0] _2409;
  wire [63:0] _2408;
  wire [63:0] _2407;
  wire [63:0] _2406;
  wire [63:0] _2405;
  wire [63:0] _2404;
  wire [63:0] _2403;
  wire [63:0] _2402;
  wire [63:0] _2401;
  wire [63:0] _2400;
  wire [63:0] _2399;
  wire [63:0] _2398;
  wire [63:0] _2397;
  wire [31:0] _2396;
  wire [63:0] _2395;
  wire [63:0] _2394;
  wire [63:0] _2393;
  wire [0:0] ifout2471;
  wire [63:0] _2392;
  wire [63:0] _2391;
  wire [63:0] _2390;
  wire [63:0] _2389;
  wire [63:0] _2388;
  wire [63:0] _2387;
  wire [7:0] _3640;
  wire [63:0] _2386;
  wire [63:0] _2385;
  wire [31:0] n_idx_3639;
  wire [31:0] _2384;
  wire [31:0] _2383;
  wire [63:0] _2382;
  wire [63:0] _2381;
  wire [63:0] _2380;
  wire [63:0] _2379;
  wire [63:0] _2378;
  wire [63:0] _2377;
  wire [63:0] _2376;
  wire [63:0] _2375;
  wire [63:0] _2374;
  wire [63:0] _2373;
  wire [63:0] _2372;
  wire [63:0] _2371;
  wire [63:0] _2370;
  wire [63:0] _2369;
  wire [63:0] _2368;
  wire [63:0] _2367;
  wire [63:0] _2366;
  wire [63:0] _2365;
  wire [63:0] _2364;
  wire [63:0] _2363;
  wire [63:0] _2362;
  wire [63:0] _2361;
  wire [63:0] _2360;
  wire [63:0] _2359;
  wire [63:0] _2358;
  wire [63:0] _2357;
  wire [63:0] _2356;
  wire [63:0] _2355;
  wire [63:0] _2354;
  wire [63:0] _2353;
  wire [63:0] _2352;
  wire [63:0] _2351;
  wire [63:0] _2350;
  wire [63:0] _2349;
  wire [63:0] _2348;
  wire [63:0] _2347;
  wire [63:0] _2346;
  wire [63:0] _2345;
  wire [63:0] _2344;
  wire [63:0] _2343;
  wire [63:0] _2342;
  wire [63:0] _2341;
  wire [63:0] _2340;
  wire [63:0] _2339;
  wire [63:0] _2338;
  wire [63:0] _2337;
  wire [63:0] _2336;
  wire [63:0] _2335;
  wire [63:0] _2334;
  wire [63:0] _2333;
  wire [63:0] _2332;
  wire [63:0] _2331;
  wire [63:0] _2330;
  wire [63:0] _2329;
  wire [63:0] _2328;
  wire [63:0] _2327;
  wire [63:0] _2326;
  wire [63:0] _2325;
  wire [63:0] _2324;
  wire [63:0] _2323;
  wire [63:0] _2322;
  wire [63:0] _2321;
  wire [63:0] _2320;
  wire [63:0] _2319;
  wire [63:0] _2318;
  wire [63:0] _2317;
  wire [63:0] _2316;
  wire [63:0] _2315;
  wire [63:0] _2314;
  wire [63:0] _2313;
  wire [63:0] _2312;
  wire [63:0] _2311;
  wire [63:0] _2310;
  wire [63:0] _2309;
  wire [63:0] _2308;
  wire [63:0] _2307;
  wire [63:0] _2306;
  wire [63:0] _2305;
  wire [63:0] _2304;
  wire [63:0] _2303;
  wire [63:0] _2302;
  wire [31:0] _2301;
  wire [63:0] _2300;
  wire [63:0] _2299;
  wire [63:0] _2298;
  wire [0:0] ifout2373;
  wire [63:0] _2297;
  wire [63:0] _2296;
  wire [63:0] _2295;
  wire [63:0] _2294;
  wire [63:0] _2293;
  wire [63:0] _2292;
  wire [7:0] _3648;
  wire [63:0] _2291;
  wire [63:0] _2290;
  wire [31:0] n_idx_3647;
  wire [31:0] _2289;
  wire [31:0] _2288;
  wire [63:0] _2287;
  wire [63:0] _2286;
  wire [63:0] _2285;
  wire [63:0] _2284;
  wire [63:0] _2283;
  wire [63:0] _2282;
  wire [63:0] _2281;
  wire [63:0] _2280;
  wire [63:0] _2279;
  wire [63:0] _2278;
  wire [63:0] _2277;
  wire [63:0] _2276;
  wire [63:0] _2275;
  wire [63:0] _2274;
  wire [63:0] _2273;
  wire [63:0] _2272;
  wire [63:0] _2271;
  wire [63:0] _2270;
  wire [63:0] _2269;
  wire [63:0] _2268;
  wire [63:0] _2267;
  wire [63:0] _2266;
  wire [63:0] _2265;
  wire [63:0] _2264;
  wire [63:0] _2263;
  wire [63:0] _2262;
  wire [63:0] _2261;
  wire [63:0] _2260;
  wire [63:0] _2259;
  wire [63:0] _2258;
  wire [63:0] _2257;
  wire [63:0] _2256;
  wire [63:0] _2255;
  wire [63:0] _2254;
  wire [63:0] _2253;
  wire [63:0] _2252;
  wire [63:0] _2251;
  wire [63:0] _2250;
  wire [63:0] _2249;
  wire [63:0] _2248;
  wire [63:0] _2247;
  wire [63:0] _2246;
  wire [63:0] _2245;
  wire [63:0] _2244;
  wire [63:0] _2243;
  wire [63:0] _2242;
  wire [63:0] _2241;
  wire [63:0] _2240;
  wire [63:0] _2239;
  wire [63:0] _2238;
  wire [63:0] _2237;
  wire [63:0] _2236;
  wire [63:0] _2235;
  wire [63:0] _2234;
  wire [63:0] _2233;
  wire [63:0] _2232;
  wire [63:0] _2231;
  wire [63:0] _2230;
  wire [63:0] _2229;
  wire [63:0] _2228;
  wire [63:0] _2227;
  wire [63:0] _2226;
  wire [63:0] _2225;
  wire [63:0] _2224;
  wire [63:0] _2223;
  wire [63:0] _2222;
  wire [63:0] _2221;
  wire [63:0] _2220;
  wire [63:0] _2219;
  wire [63:0] _2218;
  wire [63:0] _2217;
  wire [63:0] _2216;
  wire [63:0] _2215;
  wire [63:0] _2214;
  wire [63:0] _2213;
  wire [63:0] _2212;
  wire [63:0] _2211;
  wire [63:0] _2210;
  wire [63:0] _2209;
  wire [63:0] _2208;
  wire [63:0] _2207;
  wire [31:0] _2206;
  wire [63:0] _2205;
  wire [63:0] _2204;
  wire [63:0] _2203;
  wire [0:0] ifout2275;
  wire [63:0] _2202;
  wire [63:0] _2201;
  wire [63:0] _2200;
  wire [63:0] _2199;
  wire [63:0] _2198;
  wire [63:0] _2197;
  wire [7:0] _3656;
  wire [63:0] _2196;
  wire [63:0] _2195;
  wire [31:0] n_idx_3655;
  wire [31:0] _2194;
  wire [31:0] _2193;
  wire [63:0] _2192;
  wire [63:0] _2191;
  wire [63:0] _2190;
  wire [63:0] _2189;
  wire [63:0] _2188;
  wire [63:0] _2187;
  wire [63:0] _2186;
  wire [63:0] _2185;
  wire [63:0] _2184;
  wire [63:0] _2183;
  wire [63:0] _2182;
  wire [63:0] _2181;
  wire [63:0] _2180;
  wire [63:0] _2179;
  wire [63:0] _2178;
  wire [63:0] _2177;
  wire [63:0] _2176;
  wire [63:0] _2175;
  wire [63:0] _2174;
  wire [63:0] _2173;
  wire [63:0] _2172;
  wire [63:0] _2171;
  wire [63:0] _2170;
  wire [63:0] _2169;
  wire [63:0] _2168;
  wire [63:0] _2167;
  wire [63:0] _2166;
  wire [63:0] _2165;
  wire [63:0] _2164;
  wire [63:0] _2163;
  wire [63:0] _2162;
  wire [63:0] _2161;
  wire [63:0] _2160;
  wire [63:0] _2159;
  wire [63:0] _2158;
  wire [63:0] _2157;
  wire [63:0] _2156;
  wire [63:0] _2155;
  wire [63:0] _2154;
  wire [63:0] _2153;
  wire [63:0] _2152;
  wire [63:0] _2151;
  wire [63:0] _2150;
  wire [63:0] _2149;
  wire [63:0] _2148;
  wire [63:0] _2147;
  wire [63:0] _2146;
  wire [63:0] _2145;
  wire [63:0] _2144;
  wire [63:0] _2143;
  wire [63:0] _2142;
  wire [63:0] _2141;
  wire [63:0] _2140;
  wire [63:0] _2139;
  wire [63:0] _2138;
  wire [63:0] _2137;
  wire [63:0] _2136;
  wire [63:0] _2135;
  wire [63:0] _2134;
  wire [63:0] _2133;
  wire [63:0] _2132;
  wire [63:0] _2131;
  wire [63:0] _2130;
  wire [63:0] _2129;
  wire [63:0] _2128;
  wire [63:0] _2127;
  wire [63:0] _2126;
  wire [63:0] _2125;
  wire [63:0] _2124;
  wire [63:0] _2123;
  wire [63:0] _2122;
  wire [63:0] _2121;
  wire [63:0] _2120;
  wire [63:0] _2119;
  wire [63:0] _2118;
  wire [63:0] _2117;
  wire [63:0] _2116;
  wire [63:0] _2115;
  wire [63:0] _2114;
  wire [63:0] _2113;
  wire [63:0] _2112;
  wire [31:0] _2111;
  wire [63:0] _2110;
  wire [63:0] _2109;
  wire [63:0] _2108;
  wire [0:0] ifout2177;
  wire [63:0] _2107;
  wire [63:0] _2106;
  wire [63:0] _2105;
  wire [63:0] _2104;
  wire [63:0] _2103;
  wire [63:0] _2102;
  wire [7:0] _3664;
  wire [63:0] _2101;
  wire [63:0] _2100;
  wire [31:0] n_idx_3663;
  wire [31:0] _2099;
  wire [31:0] _2098;
  wire [63:0] _2097;
  wire [63:0] _2096;
  wire [63:0] _2095;
  wire [63:0] _2094;
  wire [63:0] _2093;
  wire [63:0] _2092;
  wire [63:0] _2091;
  wire [63:0] _2090;
  wire [63:0] _2089;
  wire [63:0] _2088;
  wire [63:0] _2087;
  wire [63:0] _2086;
  wire [63:0] _2085;
  wire [63:0] _2084;
  wire [63:0] _2083;
  wire [63:0] _2082;
  wire [63:0] _2081;
  wire [63:0] _2080;
  wire [63:0] _2079;
  wire [63:0] _2078;
  wire [63:0] _2077;
  wire [63:0] _2076;
  wire [63:0] _2075;
  wire [63:0] _2074;
  wire [63:0] _2073;
  wire [63:0] _2072;
  wire [63:0] _2071;
  wire [63:0] _2070;
  wire [63:0] _2069;
  wire [63:0] _2068;
  wire [63:0] _2067;
  wire [63:0] _2066;
  wire [63:0] _2065;
  wire [63:0] _2064;
  wire [63:0] _2063;
  wire [63:0] _2062;
  wire [63:0] _2061;
  wire [63:0] _2060;
  wire [63:0] _2059;
  wire [63:0] _2058;
  wire [63:0] _2057;
  wire [63:0] _2056;
  wire [63:0] _2055;
  wire [63:0] _2054;
  wire [63:0] _2053;
  wire [63:0] _2052;
  wire [63:0] _2051;
  wire [63:0] _2050;
  wire [63:0] _2049;
  wire [63:0] _2048;
  wire [63:0] _2047;
  wire [63:0] _2046;
  wire [63:0] _2045;
  wire [63:0] _2044;
  wire [63:0] _2043;
  wire [63:0] _2042;
  wire [63:0] _2041;
  wire [63:0] _2040;
  wire [63:0] _2039;
  wire [63:0] _2038;
  wire [63:0] _2037;
  wire [63:0] _2036;
  wire [63:0] _2035;
  wire [63:0] _2034;
  wire [63:0] _2033;
  wire [63:0] _2032;
  wire [63:0] _2031;
  wire [63:0] _2030;
  wire [63:0] _2029;
  wire [63:0] _2028;
  wire [63:0] _2027;
  wire [63:0] _2026;
  wire [63:0] _2025;
  wire [63:0] _2024;
  wire [63:0] _2023;
  wire [63:0] _2022;
  wire [63:0] _2021;
  wire [63:0] _2020;
  wire [63:0] _2019;
  wire [63:0] _2018;
  wire [63:0] _2017;
  wire [31:0] _2016;
  wire [63:0] _2015;
  wire [63:0] _2014;
  wire [63:0] _2013;
  wire [0:0] ifout2079;
  wire [63:0] _2012;
  wire [63:0] _2011;
  wire [63:0] _2010;
  wire [63:0] _2009;
  wire [63:0] _2008;
  wire [63:0] _2007;
  wire [7:0] _3672;
  wire [63:0] _2006;
  wire [63:0] _2005;
  wire [31:0] n_idx_3671;
  wire [31:0] _2004;
  wire [31:0] _2003;
  wire [63:0] _2002;
  wire [63:0] _2001;
  wire [63:0] _2000;
  wire [63:0] _1999;
  wire [63:0] _1998;
  wire [63:0] _1997;
  wire [63:0] _1996;
  wire [63:0] _1995;
  wire [63:0] _1994;
  wire [63:0] _1993;
  wire [63:0] _1992;
  wire [63:0] _1991;
  wire [63:0] _1990;
  wire [63:0] _1989;
  wire [63:0] _1988;
  wire [63:0] _1987;
  wire [63:0] _1986;
  wire [63:0] _1985;
  wire [63:0] _1984;
  wire [63:0] _1983;
  wire [63:0] _1982;
  wire [63:0] _1981;
  wire [63:0] _1980;
  wire [63:0] _1979;
  wire [63:0] _1978;
  wire [63:0] _1977;
  wire [63:0] _1976;
  wire [63:0] _1975;
  wire [63:0] _1974;
  wire [63:0] _1973;
  wire [63:0] _1972;
  wire [63:0] _1971;
  wire [63:0] _1970;
  wire [63:0] _1969;
  wire [63:0] _1968;
  wire [63:0] _1967;
  wire [63:0] _1966;
  wire [63:0] _1965;
  wire [63:0] _1964;
  wire [63:0] _1963;
  wire [63:0] _1962;
  wire [63:0] _1961;
  wire [63:0] _1960;
  wire [63:0] _1959;
  wire [63:0] _1958;
  wire [63:0] _1957;
  wire [63:0] _1956;
  wire [63:0] _1955;
  wire [63:0] _1954;
  wire [63:0] _1953;
  wire [63:0] _1952;
  wire [63:0] _1951;
  wire [63:0] _1950;
  wire [63:0] _1949;
  wire [63:0] _1948;
  wire [63:0] _1947;
  wire [63:0] _1946;
  wire [63:0] _1945;
  wire [63:0] _1944;
  wire [63:0] _1943;
  wire [63:0] _1942;
  wire [63:0] _1941;
  wire [63:0] _1940;
  wire [63:0] _1939;
  wire [63:0] _1938;
  wire [63:0] _1937;
  wire [63:0] _1936;
  wire [63:0] _1935;
  wire [63:0] _1934;
  wire [63:0] _1933;
  wire [63:0] _1932;
  wire [63:0] _1931;
  wire [63:0] _1930;
  wire [63:0] _1929;
  wire [63:0] _1928;
  wire [63:0] _1927;
  wire [63:0] _1926;
  wire [63:0] _1925;
  wire [63:0] _1924;
  wire [63:0] _1923;
  wire [63:0] _1922;
  wire [31:0] _1921;
  wire [63:0] _1920;
  wire [63:0] _1919;
  wire [63:0] _1918;
  wire [0:0] ifout1981;
  wire [63:0] _1917;
  wire [63:0] _1916;
  wire [63:0] _1915;
  wire [63:0] _1914;
  wire [63:0] _1913;
  wire [63:0] _1912;
  wire [7:0] _3680;
  wire [63:0] _1911;
  wire [63:0] _1910;
  wire [31:0] n_idx_3679;
  wire [31:0] _1909;
  wire [31:0] _1908;
  wire [63:0] _1907;
  wire [63:0] _1906;
  wire [63:0] _1905;
  wire [63:0] _1904;
  wire [63:0] _1903;
  wire [63:0] _1902;
  wire [63:0] _1901;
  wire [63:0] _1900;
  wire [63:0] _1899;
  wire [63:0] _1898;
  wire [63:0] _1897;
  wire [63:0] _1896;
  wire [63:0] _1895;
  wire [63:0] _1894;
  wire [63:0] _1893;
  wire [63:0] _1892;
  wire [63:0] _1891;
  wire [63:0] _1890;
  wire [63:0] _1889;
  wire [63:0] _1888;
  wire [63:0] _1887;
  wire [63:0] _1886;
  wire [63:0] _1885;
  wire [63:0] _1884;
  wire [63:0] _1883;
  wire [63:0] _1882;
  wire [63:0] _1881;
  wire [63:0] _1880;
  wire [63:0] _1879;
  wire [63:0] _1878;
  wire [63:0] _1877;
  wire [63:0] _1876;
  wire [63:0] _1875;
  wire [63:0] _1874;
  wire [63:0] _1873;
  wire [63:0] _1872;
  wire [63:0] _1871;
  wire [63:0] _1870;
  wire [63:0] _1869;
  wire [63:0] _1868;
  wire [63:0] _1867;
  wire [63:0] _1866;
  wire [63:0] _1865;
  wire [63:0] _1864;
  wire [63:0] _1863;
  wire [63:0] _1862;
  wire [63:0] _1861;
  wire [63:0] _1860;
  wire [63:0] _1859;
  wire [63:0] _1858;
  wire [63:0] _1857;
  wire [63:0] _1856;
  wire [63:0] _1855;
  wire [63:0] _1854;
  wire [63:0] _1853;
  wire [63:0] _1852;
  wire [63:0] _1851;
  wire [63:0] _1850;
  wire [63:0] _1849;
  wire [63:0] _1848;
  wire [63:0] _1847;
  wire [63:0] _1846;
  wire [63:0] _1845;
  wire [63:0] _1844;
  wire [63:0] _1843;
  wire [63:0] _1842;
  wire [63:0] _1841;
  wire [63:0] _1840;
  wire [63:0] _1839;
  wire [63:0] _1838;
  wire [63:0] _1837;
  wire [63:0] _1836;
  wire [63:0] _1835;
  wire [63:0] _1834;
  wire [63:0] _1833;
  wire [63:0] _1832;
  wire [63:0] _1831;
  wire [63:0] _1830;
  wire [63:0] _1829;
  wire [63:0] _1828;
  wire [63:0] _1827;
  wire [31:0] _1826;
  wire [63:0] _1825;
  wire [63:0] _1824;
  wire [63:0] _1823;
  wire [0:0] ifout1883;
  wire [63:0] _1822;
  wire [63:0] _1821;
  wire [63:0] _1820;
  wire [63:0] _1819;
  wire [63:0] _1818;
  wire [63:0] _1817;
  wire [7:0] _3687;
  wire [63:0] _1816;
  wire [63:0] _1815;
  wire [31:0] n_idx_3686;
  wire [31:0] _1814;
  wire [31:0] _1813;
  wire [63:0] _1812;
  wire [63:0] _1811;
  wire [63:0] _1810;
  wire [63:0] _1809;
  wire [63:0] _1808;
  wire [63:0] _1807;
  wire [63:0] _1806;
  wire [63:0] _1805;
  wire [63:0] _1804;
  wire [63:0] _1803;
  wire [63:0] _1802;
  wire [63:0] _1801;
  wire [63:0] _1800;
  wire [63:0] _1799;
  wire [63:0] _1798;
  wire [63:0] _1797;
  wire [63:0] _1796;
  wire [63:0] _1795;
  wire [63:0] _1794;
  wire [63:0] _1793;
  wire [63:0] _1792;
  wire [63:0] _1791;
  wire [63:0] _1790;
  wire [63:0] _1789;
  wire [63:0] _1788;
  wire [63:0] _1787;
  wire [63:0] _1786;
  wire [63:0] _1785;
  wire [63:0] _1784;
  wire [63:0] _1783;
  wire [63:0] _1782;
  wire [63:0] _1781;
  wire [63:0] _1780;
  wire [63:0] _1779;
  wire [63:0] _1778;
  wire [63:0] _1777;
  wire [63:0] _1776;
  wire [63:0] _1775;
  wire [63:0] _1774;
  wire [63:0] _1773;
  wire [63:0] _1772;
  wire [63:0] _1771;
  wire [63:0] _1770;
  wire [63:0] _1769;
  wire [63:0] _1768;
  wire [63:0] _1767;
  wire [63:0] _1766;
  wire [63:0] _1765;
  wire [63:0] _1764;
  wire [63:0] _1763;
  wire [63:0] _1762;
  wire [63:0] _1761;
  wire [63:0] _1760;
  wire [63:0] _1759;
  wire [63:0] _1758;
  wire [63:0] _1757;
  wire [63:0] _1756;
  wire [63:0] _1755;
  wire [63:0] _1754;
  wire [63:0] _1753;
  wire [63:0] _1752;
  wire [63:0] _1751;
  wire [63:0] _1750;
  wire [63:0] _1749;
  wire [63:0] _1748;
  wire [63:0] _1747;
  wire [63:0] _1746;
  wire [63:0] _1745;
  wire [63:0] _1744;
  wire [63:0] _1743;
  wire [63:0] _1742;
  wire [63:0] _1741;
  wire [63:0] _1740;
  wire [63:0] _1739;
  wire [63:0] _1738;
  wire [63:0] _1737;
  wire [63:0] _1736;
  wire [63:0] _1735;
  wire [63:0] _1734;
  wire [63:0] _1733;
  wire [63:0] _1732;
  wire [31:0] _1731;
  wire [63:0] _1730;
  wire [63:0] _1729;
  wire [63:0] _1728;
  wire [0:0] ifout1785;
  wire [63:0] _1727;
  wire [63:0] _1726;
  wire [63:0] _1725;
  wire [63:0] _1724;
  wire [63:0] _1723;
  wire [63:0] _1722;
  wire [31:0] off_3683;
  wire [31:0] _1721;
  wire [63:0] _1720;
  wire [31:0] idx_3682;
  wire [31:0] _1719;
  wire [31:0] _1718;
  wire [63:0] _1717;
  wire [63:0] _1716;
  wire [63:0] _1715;
  wire [63:0] _1714;
  wire [63:0] _1713;
  wire [63:0] _1712;
  wire [63:0] _1711;
  wire [63:0] _1710;
  wire [63:0] _1709;
  wire [63:0] _1708;
  wire [63:0] _1707;
  wire [63:0] _1706;
  wire [63:0] _1705;
  wire [63:0] _1704;
  wire [63:0] _1703;
  wire [63:0] _1702;
  wire [63:0] _1701;
  wire [63:0] _1700;
  wire [63:0] _1699;
  wire [63:0] _1698;
  wire [63:0] _1697;
  wire [63:0] _1696;
  wire [63:0] _1695;
  wire [63:0] _1694;
  wire [63:0] _1693;
  wire [63:0] _1692;
  wire [63:0] _1691;
  wire [63:0] _1690;
  wire [63:0] _1689;
  wire [63:0] _1688;
  wire [63:0] _1687;
  wire [63:0] _1686;
  wire [63:0] _1685;
  wire [63:0] _1684;
  wire [63:0] _1683;
  wire [63:0] _1682;
  wire [63:0] _1681;
  wire [63:0] _1680;
  wire [63:0] _1679;
  wire [63:0] _1678;
  wire [63:0] _1677;
  wire [63:0] _1676;
  wire [63:0] _1675;
  wire [63:0] _1674;
  wire [63:0] _1673;
  wire [63:0] _1672;
  wire [63:0] _1671;
  wire [63:0] _1670;
  wire [63:0] _1669;
  wire [63:0] _1668;
  wire [63:0] _1667;
  wire [63:0] _1666;
  wire [63:0] _1665;
  wire [63:0] _1664;
  wire [63:0] _1663;
  wire [63:0] _1662;
  wire [63:0] _1661;
  wire [63:0] _1660;
  wire [63:0] _1659;
  wire [63:0] _1658;
  wire [63:0] _1657;
  wire [63:0] _1656;
  wire [63:0] _1655;
  wire [63:0] _1654;
  wire [63:0] _1653;
  wire [63:0] _1652;
  wire [63:0] _1651;
  wire [63:0] _1650;
  wire [63:0] _1649;
  wire [63:0] _1648;
  wire [63:0] _1647;
  wire [63:0] _1646;
  wire [63:0] _1645;
  wire [63:0] _1644;
  wire [63:0] _1643;
  wire [63:0] _1642;
  wire [63:0] _1641;
  wire [63:0] _1640;
  wire [63:0] _1639;
  wire [63:0] _1638;
  wire [63:0] _1637;
  wire [31:0] _1636;
  wire [63:0] _1635;
  wire [63:0] _1634;
  wire [63:0] _1633;
  wire [0:0] ifout1687;
  wire [63:0] _1632;
  wire [63:0] _1631;
  wire [63:0] _1630;
  wire [63:0] _1629;
  wire [63:0] _1628;
  wire [63:0] _1627;
  wire [31:0] off_3675;
  wire [31:0] _1626;
  wire [63:0] _1625;
  wire [31:0] idx_3674;
  wire [31:0] _1624;
  wire [31:0] _1623;
  wire [63:0] _1622;
  wire [63:0] _1621;
  wire [63:0] _1620;
  wire [63:0] _1619;
  wire [63:0] _1618;
  wire [63:0] _1617;
  wire [63:0] _1616;
  wire [63:0] _1615;
  wire [63:0] _1614;
  wire [63:0] _1613;
  wire [63:0] _1612;
  wire [63:0] _1611;
  wire [63:0] _1610;
  wire [63:0] _1609;
  wire [63:0] _1608;
  wire [63:0] _1607;
  wire [63:0] _1606;
  wire [63:0] _1605;
  wire [63:0] _1604;
  wire [63:0] _1603;
  wire [63:0] _1602;
  wire [63:0] _1601;
  wire [63:0] _1600;
  wire [63:0] _1599;
  wire [63:0] _1598;
  wire [63:0] _1597;
  wire [63:0] _1596;
  wire [63:0] _1595;
  wire [63:0] _1594;
  wire [63:0] _1593;
  wire [63:0] _1592;
  wire [63:0] _1591;
  wire [63:0] _1590;
  wire [63:0] _1589;
  wire [63:0] _1588;
  wire [63:0] _1587;
  wire [63:0] _1586;
  wire [63:0] _1585;
  wire [63:0] _1584;
  wire [63:0] _1583;
  wire [63:0] _1582;
  wire [63:0] _1581;
  wire [63:0] _1580;
  wire [63:0] _1579;
  wire [63:0] _1578;
  wire [63:0] _1577;
  wire [63:0] _1576;
  wire [63:0] _1575;
  wire [63:0] _1574;
  wire [63:0] _1573;
  wire [63:0] _1572;
  wire [63:0] _1571;
  wire [63:0] _1570;
  wire [63:0] _1569;
  wire [63:0] _1568;
  wire [63:0] _1567;
  wire [63:0] _1566;
  wire [63:0] _1565;
  wire [63:0] _1564;
  wire [63:0] _1563;
  wire [63:0] _1562;
  wire [63:0] _1561;
  wire [63:0] _1560;
  wire [63:0] _1559;
  wire [63:0] _1558;
  wire [63:0] _1557;
  wire [63:0] _1556;
  wire [63:0] _1555;
  wire [63:0] _1554;
  wire [63:0] _1553;
  wire [63:0] _1552;
  wire [63:0] _1551;
  wire [63:0] _1550;
  wire [63:0] _1549;
  wire [63:0] _1548;
  wire [63:0] _1547;
  wire [63:0] _1546;
  wire [63:0] _1545;
  wire [63:0] _1544;
  wire [63:0] _1543;
  wire [63:0] _1542;
  wire [31:0] _1541;
  wire [63:0] _1540;
  wire [63:0] _1539;
  wire [63:0] _1538;
  wire [0:0] ifout1589;
  wire [63:0] _1537;
  wire [63:0] _1536;
  wire [63:0] _1535;
  wire [63:0] _1534;
  wire [63:0] _1533;
  wire [63:0] _1532;
  wire [31:0] off_3667;
  wire [31:0] _1531;
  wire [63:0] _1530;
  wire [31:0] idx_3666;
  wire [31:0] _1529;
  wire [31:0] _1528;
  wire [63:0] _1527;
  wire [63:0] _1526;
  wire [63:0] _1525;
  wire [63:0] _1524;
  wire [63:0] _1523;
  wire [63:0] _1522;
  wire [63:0] _1521;
  wire [63:0] _1520;
  wire [63:0] _1519;
  wire [63:0] _1518;
  wire [63:0] _1517;
  wire [63:0] _1516;
  wire [63:0] _1515;
  wire [63:0] _1514;
  wire [63:0] _1513;
  wire [63:0] _1512;
  wire [63:0] _1511;
  wire [63:0] _1510;
  wire [63:0] _1509;
  wire [63:0] _1508;
  wire [63:0] _1507;
  wire [63:0] _1506;
  wire [63:0] _1505;
  wire [63:0] _1504;
  wire [63:0] _1503;
  wire [63:0] _1502;
  wire [63:0] _1501;
  wire [63:0] _1500;
  wire [63:0] _1499;
  wire [63:0] _1498;
  wire [63:0] _1497;
  wire [63:0] _1496;
  wire [63:0] _1495;
  wire [63:0] _1494;
  wire [63:0] _1493;
  wire [63:0] _1492;
  wire [63:0] _1491;
  wire [63:0] _1490;
  wire [63:0] _1489;
  wire [63:0] _1488;
  wire [63:0] _1487;
  wire [63:0] _1486;
  wire [63:0] _1485;
  wire [63:0] _1484;
  wire [63:0] _1483;
  wire [63:0] _1482;
  wire [63:0] _1481;
  wire [63:0] _1480;
  wire [63:0] _1479;
  wire [63:0] _1478;
  wire [63:0] _1477;
  wire [63:0] _1476;
  wire [63:0] _1475;
  wire [63:0] _1474;
  wire [63:0] _1473;
  wire [63:0] _1472;
  wire [63:0] _1471;
  wire [63:0] _1470;
  wire [63:0] _1469;
  wire [63:0] _1468;
  wire [63:0] _1467;
  wire [63:0] _1466;
  wire [63:0] _1465;
  wire [63:0] _1464;
  wire [63:0] _1463;
  wire [63:0] _1462;
  wire [63:0] _1461;
  wire [63:0] _1460;
  wire [63:0] _1459;
  wire [63:0] _1458;
  wire [63:0] _1457;
  wire [63:0] _1456;
  wire [63:0] _1455;
  wire [63:0] _1454;
  wire [63:0] _1453;
  wire [63:0] _1452;
  wire [63:0] _1451;
  wire [63:0] _1450;
  wire [63:0] _1449;
  wire [63:0] _1448;
  wire [63:0] _1447;
  wire [31:0] _1446;
  wire [63:0] _1445;
  wire [63:0] _1444;
  wire [63:0] _1443;
  wire [0:0] ifout1491;
  wire [63:0] _1442;
  wire [63:0] _1441;
  wire [63:0] _1440;
  wire [63:0] _1439;
  wire [63:0] _1438;
  wire [63:0] _1437;
  wire [31:0] off_3659;
  wire [31:0] _1436;
  wire [63:0] _1435;
  wire [31:0] idx_3658;
  wire [31:0] _1434;
  wire [31:0] _1433;
  wire [63:0] _1432;
  wire [63:0] _1431;
  wire [63:0] _1430;
  wire [63:0] _1429;
  wire [63:0] _1428;
  wire [63:0] _1427;
  wire [63:0] _1426;
  wire [63:0] _1425;
  wire [63:0] _1424;
  wire [63:0] _1423;
  wire [63:0] _1422;
  wire [63:0] _1421;
  wire [63:0] _1420;
  wire [63:0] _1419;
  wire [63:0] _1418;
  wire [63:0] _1417;
  wire [63:0] _1416;
  wire [63:0] _1415;
  wire [63:0] _1414;
  wire [63:0] _1413;
  wire [63:0] _1412;
  wire [63:0] _1411;
  wire [63:0] _1410;
  wire [63:0] _1409;
  wire [63:0] _1408;
  wire [63:0] _1407;
  wire [63:0] _1406;
  wire [63:0] _1405;
  wire [63:0] _1404;
  wire [63:0] _1403;
  wire [63:0] _1402;
  wire [63:0] _1401;
  wire [63:0] _1400;
  wire [63:0] _1399;
  wire [63:0] _1398;
  wire [63:0] _1397;
  wire [63:0] _1396;
  wire [63:0] _1395;
  wire [63:0] _1394;
  wire [63:0] _1393;
  wire [63:0] _1392;
  wire [63:0] _1391;
  wire [63:0] _1390;
  wire [63:0] _1389;
  wire [63:0] _1388;
  wire [63:0] _1387;
  wire [63:0] _1386;
  wire [63:0] _1385;
  wire [63:0] _1384;
  wire [63:0] _1383;
  wire [63:0] _1382;
  wire [63:0] _1381;
  wire [63:0] _1380;
  wire [63:0] _1379;
  wire [63:0] _1378;
  wire [63:0] _1377;
  wire [63:0] _1376;
  wire [63:0] _1375;
  wire [63:0] _1374;
  wire [63:0] _1373;
  wire [63:0] _1372;
  wire [63:0] _1371;
  wire [63:0] _1370;
  wire [63:0] _1369;
  wire [63:0] _1368;
  wire [63:0] _1367;
  wire [63:0] _1366;
  wire [63:0] _1365;
  wire [63:0] _1364;
  wire [63:0] _1363;
  wire [63:0] _1362;
  wire [63:0] _1361;
  wire [63:0] _1360;
  wire [63:0] _1359;
  wire [63:0] _1358;
  wire [63:0] _1357;
  wire [63:0] _1356;
  wire [63:0] _1355;
  wire [63:0] _1354;
  wire [63:0] _1353;
  wire [63:0] _1352;
  wire [31:0] _1351;
  wire [63:0] _1350;
  wire [63:0] _1349;
  wire [63:0] _1348;
  wire [0:0] ifout1393;
  wire [63:0] _1347;
  wire [63:0] _1346;
  wire [63:0] _1345;
  wire [63:0] _1344;
  wire [63:0] _1343;
  wire [63:0] _1342;
  wire [31:0] off_3651;
  wire [31:0] _1341;
  wire [63:0] _1340;
  wire [31:0] idx_3650;
  wire [31:0] _1339;
  wire [31:0] _1338;
  wire [63:0] _1337;
  wire [63:0] _1336;
  wire [63:0] _1335;
  wire [63:0] _1334;
  wire [63:0] _1333;
  wire [63:0] _1332;
  wire [63:0] _1331;
  wire [63:0] _1330;
  wire [63:0] _1329;
  wire [63:0] _1328;
  wire [63:0] _1327;
  wire [63:0] _1326;
  wire [63:0] _1325;
  wire [63:0] _1324;
  wire [63:0] _1323;
  wire [63:0] _1322;
  wire [63:0] _1321;
  wire [63:0] _1320;
  wire [63:0] _1319;
  wire [63:0] _1318;
  wire [63:0] _1317;
  wire [63:0] _1316;
  wire [63:0] _1315;
  wire [63:0] _1314;
  wire [63:0] _1313;
  wire [63:0] _1312;
  wire [63:0] _1311;
  wire [63:0] _1310;
  wire [63:0] _1309;
  wire [63:0] _1308;
  wire [63:0] _1307;
  wire [63:0] _1306;
  wire [63:0] _1305;
  wire [63:0] _1304;
  wire [63:0] _1303;
  wire [63:0] _1302;
  wire [63:0] _1301;
  wire [63:0] _1300;
  wire [63:0] _1299;
  wire [63:0] _1298;
  wire [63:0] _1297;
  wire [63:0] _1296;
  wire [63:0] _1295;
  wire [63:0] _1294;
  wire [63:0] _1293;
  wire [63:0] _1292;
  wire [63:0] _1291;
  wire [63:0] _1290;
  wire [63:0] _1289;
  wire [63:0] _1288;
  wire [63:0] _1287;
  wire [63:0] _1286;
  wire [63:0] _1285;
  wire [63:0] _1284;
  wire [63:0] _1283;
  wire [63:0] _1282;
  wire [63:0] _1281;
  wire [63:0] _1280;
  wire [63:0] _1279;
  wire [63:0] _1278;
  wire [63:0] _1277;
  wire [63:0] _1276;
  wire [63:0] _1275;
  wire [63:0] _1274;
  wire [63:0] _1273;
  wire [63:0] _1272;
  wire [63:0] _1271;
  wire [63:0] _1270;
  wire [63:0] _1269;
  wire [63:0] _1268;
  wire [63:0] _1267;
  wire [63:0] _1266;
  wire [63:0] _1265;
  wire [63:0] _1264;
  wire [63:0] _1263;
  wire [63:0] _1262;
  wire [63:0] _1261;
  wire [63:0] _1260;
  wire [63:0] _1259;
  wire [63:0] _1258;
  wire [63:0] _1257;
  wire [31:0] _1256;
  wire [63:0] _1255;
  wire [63:0] _1254;
  wire [63:0] _1253;
  wire [0:0] ifout1295;
  wire [63:0] _1252;
  wire [63:0] _1251;
  wire [63:0] _1250;
  wire [63:0] _1249;
  wire [63:0] _1248;
  wire [63:0] _1247;
  wire [31:0] off_3643;
  wire [31:0] _1246;
  wire [63:0] _1245;
  wire [31:0] idx_3642;
  wire [31:0] _1244;
  wire [31:0] _1243;
  wire [63:0] _1242;
  wire [63:0] _1241;
  wire [63:0] _1240;
  wire [63:0] _1239;
  wire [63:0] _1238;
  wire [63:0] _1237;
  wire [63:0] _1236;
  wire [63:0] _1235;
  wire [63:0] _1234;
  wire [63:0] _1233;
  wire [63:0] _1232;
  wire [63:0] _1231;
  wire [63:0] _1230;
  wire [63:0] _1229;
  wire [63:0] _1228;
  wire [63:0] _1227;
  wire [63:0] _1226;
  wire [63:0] _1225;
  wire [63:0] _1224;
  wire [63:0] _1223;
  wire [63:0] _1222;
  wire [63:0] _1221;
  wire [63:0] _1220;
  wire [63:0] _1219;
  wire [63:0] _1218;
  wire [63:0] _1217;
  wire [63:0] _1216;
  wire [63:0] _1215;
  wire [63:0] _1214;
  wire [63:0] _1213;
  wire [63:0] _1212;
  wire [63:0] _1211;
  wire [63:0] _1210;
  wire [63:0] _1209;
  wire [63:0] _1208;
  wire [63:0] _1207;
  wire [63:0] _1206;
  wire [63:0] _1205;
  wire [63:0] _1204;
  wire [63:0] _1203;
  wire [63:0] _1202;
  wire [63:0] _1201;
  wire [63:0] _1200;
  wire [63:0] _1199;
  wire [63:0] _1198;
  wire [63:0] _1197;
  wire [63:0] _1196;
  wire [63:0] _1195;
  wire [63:0] _1194;
  wire [63:0] _1193;
  wire [63:0] _1192;
  wire [63:0] _1191;
  wire [63:0] _1190;
  wire [63:0] _1189;
  wire [63:0] _1188;
  wire [63:0] _1187;
  wire [63:0] _1186;
  wire [63:0] _1185;
  wire [63:0] _1184;
  wire [63:0] _1183;
  wire [63:0] _1182;
  wire [63:0] _1181;
  wire [63:0] _1180;
  wire [63:0] _1179;
  wire [63:0] _1178;
  wire [63:0] _1177;
  wire [63:0] _1176;
  wire [63:0] _1175;
  wire [63:0] _1174;
  wire [63:0] _1173;
  wire [63:0] _1172;
  wire [63:0] _1171;
  wire [63:0] _1170;
  wire [63:0] _1169;
  wire [63:0] _1168;
  wire [63:0] _1167;
  wire [63:0] _1166;
  wire [63:0] _1165;
  wire [63:0] _1164;
  wire [63:0] _1163;
  wire [63:0] _1162;
  wire [31:0] _1161;
  wire [63:0] _1160;
  wire [63:0] _1159;
  wire [63:0] _1158;
  wire [0:0] ifout1197;
  wire [63:0] _1157;
  wire [63:0] _1156;
  wire [63:0] _1155;
  wire [63:0] _1154;
  wire [63:0] _1153;
  wire [63:0] _1152;
  wire [31:0] off_3635;
  wire [31:0] _1151;
  wire [63:0] _1150;
  wire [31:0] idx_3634;
  wire [31:0] _1149;
  wire [31:0] _1148;
  wire [63:0] _1147;
  wire [63:0] _1146;
  wire [63:0] _1145;
  wire [63:0] _1144;
  wire [63:0] _1143;
  wire [63:0] _1142;
  wire [63:0] _1141;
  wire [63:0] _1140;
  wire [63:0] _1139;
  wire [63:0] _1138;
  wire [63:0] _1137;
  wire [63:0] _1136;
  wire [63:0] _1135;
  wire [63:0] _1134;
  wire [63:0] _1133;
  wire [63:0] _1132;
  wire [63:0] _1131;
  wire [63:0] _1130;
  wire [63:0] _1129;
  wire [63:0] _1128;
  wire [63:0] _1127;
  wire [63:0] _1126;
  wire [63:0] _1125;
  wire [63:0] _1124;
  wire [63:0] _1123;
  wire [63:0] _1122;
  wire [63:0] _1121;
  wire [63:0] _1120;
  wire [63:0] _1119;
  wire [63:0] _1118;
  wire [63:0] _1117;
  wire [63:0] _1116;
  wire [63:0] _1115;
  wire [63:0] _1114;
  wire [63:0] _1113;
  wire [63:0] _1112;
  wire [63:0] _1111;
  wire [63:0] _1110;
  wire [63:0] _1109;
  wire [63:0] _1108;
  wire [63:0] _1107;
  wire [63:0] _1106;
  wire [63:0] _1105;
  wire [63:0] _1104;
  wire [63:0] _1103;
  wire [63:0] _1102;
  wire [63:0] _1101;
  wire [63:0] _1100;
  wire [63:0] _1099;
  wire [63:0] _1098;
  wire [63:0] _1097;
  wire [63:0] _1096;
  wire [63:0] _1095;
  wire [63:0] _1094;
  wire [63:0] _1093;
  wire [63:0] _1092;
  wire [63:0] _1091;
  wire [63:0] _1090;
  wire [63:0] _1089;
  wire [63:0] _1088;
  wire [63:0] _1087;
  wire [63:0] _1086;
  wire [63:0] _1085;
  wire [63:0] _1084;
  wire [63:0] _1083;
  wire [63:0] _1082;
  wire [63:0] _1081;
  wire [63:0] _1080;
  wire [63:0] _1079;
  wire [63:0] _1078;
  wire [63:0] _1077;
  wire [63:0] _1076;
  wire [63:0] _1075;
  wire [63:0] _1074;
  wire [63:0] _1073;
  wire [63:0] _1072;
  wire [63:0] _1071;
  wire [63:0] _1070;
  wire [63:0] _1069;
  wire [63:0] _1068;
  wire [63:0] _1067;
  wire [31:0] _1066;
  wire [63:0] _1065;
  wire [63:0] _1064;
  wire [63:0] _1063;
  wire [0:0] ifout1099;
  wire [63:0] _1062;
  wire [63:0] _1061;
  wire [63:0] _1060;
  wire [63:0] _1059;
  wire [63:0] _1058;
  wire [63:0] _1057;
  wire [31:0] off_3627;
  wire [31:0] _1056;
  wire [63:0] _1055;
  wire [31:0] idx_3626;
  wire [31:0] _1054;
  wire [31:0] _1053;
  wire [63:0] _1052;
  wire [63:0] _1051;
  wire [63:0] _1050;
  wire [63:0] _1049;
  wire [63:0] _1048;
  wire [63:0] _1047;
  wire [63:0] _1046;
  wire [63:0] _1045;
  wire [63:0] _1044;
  wire [63:0] _1043;
  wire [63:0] _1042;
  wire [63:0] _1041;
  wire [63:0] _1040;
  wire [63:0] _1039;
  wire [63:0] _1038;
  wire [63:0] _1037;
  wire [63:0] _1036;
  wire [63:0] _1035;
  wire [63:0] _1034;
  wire [63:0] _1033;
  wire [63:0] _1032;
  wire [63:0] _1031;
  wire [63:0] _1030;
  wire [63:0] _1029;
  wire [63:0] _1028;
  wire [63:0] _1027;
  wire [63:0] _1026;
  wire [63:0] _1025;
  wire [63:0] _1024;
  wire [63:0] _1023;
  wire [63:0] _1022;
  wire [63:0] _1021;
  wire [63:0] _1020;
  wire [63:0] _1019;
  wire [63:0] _1018;
  wire [63:0] _1017;
  wire [63:0] _1016;
  wire [63:0] _1015;
  wire [63:0] _1014;
  wire [63:0] _1013;
  wire [63:0] _1012;
  wire [63:0] _1011;
  wire [63:0] _1010;
  wire [63:0] _1009;
  wire [63:0] _1008;
  wire [63:0] _1007;
  wire [63:0] _1006;
  wire [63:0] _1005;
  wire [63:0] _1004;
  wire [63:0] _1003;
  wire [63:0] _1002;
  wire [63:0] _1001;
  wire [63:0] _1000;
  wire [63:0] _999;
  wire [63:0] _998;
  wire [63:0] _997;
  wire [63:0] _996;
  wire [63:0] _995;
  wire [63:0] _994;
  wire [63:0] _993;
  wire [63:0] _992;
  wire [63:0] _991;
  wire [63:0] _990;
  wire [63:0] _989;
  wire [63:0] _988;
  wire [63:0] _987;
  wire [63:0] _986;
  wire [63:0] _985;
  wire [63:0] _984;
  wire [63:0] _983;
  wire [63:0] _982;
  wire [63:0] _981;
  wire [63:0] _980;
  wire [63:0] _979;
  wire [63:0] _978;
  wire [63:0] _977;
  wire [63:0] _976;
  wire [63:0] _975;
  wire [63:0] _974;
  wire [63:0] _973;
  wire [63:0] _972;
  wire [31:0] _971;
  wire [63:0] _970;
  wire [63:0] _969;
  wire [63:0] _968;
  wire [0:0] ifout1001;
  wire [63:0] _967;
  wire [63:0] _966;
  wire [63:0] _965;
  wire [63:0] _964;
  wire [63:0] _963;
  wire [63:0] _962;
  wire [31:0] off_3619;
  wire [31:0] _961;
  wire [63:0] _960;
  wire [31:0] idx_3618;
  wire [31:0] _959;
  wire [31:0] _958;
  wire [63:0] _957;
  wire [63:0] _956;
  wire [63:0] _955;
  wire [63:0] _954;
  wire [63:0] _953;
  wire [63:0] _952;
  wire [63:0] _951;
  wire [63:0] _950;
  wire [63:0] _949;
  wire [63:0] _948;
  wire [63:0] _947;
  wire [63:0] _946;
  wire [63:0] _945;
  wire [63:0] _944;
  wire [63:0] _943;
  wire [63:0] _942;
  wire [63:0] _941;
  wire [63:0] _940;
  wire [63:0] _939;
  wire [63:0] _938;
  wire [63:0] _937;
  wire [63:0] _936;
  wire [63:0] _935;
  wire [63:0] _934;
  wire [63:0] _933;
  wire [63:0] _932;
  wire [63:0] _931;
  wire [63:0] _930;
  wire [63:0] _929;
  wire [63:0] _928;
  wire [63:0] _927;
  wire [63:0] _926;
  wire [63:0] _925;
  wire [63:0] _924;
  wire [63:0] _923;
  wire [63:0] _922;
  wire [63:0] _921;
  wire [63:0] _920;
  wire [63:0] _919;
  wire [63:0] _918;
  wire [63:0] _917;
  wire [63:0] _916;
  wire [63:0] _915;
  wire [63:0] _914;
  wire [63:0] _913;
  wire [63:0] _912;
  wire [63:0] _911;
  wire [63:0] _910;
  wire [63:0] _909;
  wire [63:0] _908;
  wire [63:0] _907;
  wire [63:0] _906;
  wire [63:0] _905;
  wire [63:0] _904;
  wire [63:0] _903;
  wire [63:0] _902;
  wire [63:0] _901;
  wire [63:0] _900;
  wire [63:0] _899;
  wire [63:0] _898;
  wire [63:0] _897;
  wire [63:0] _896;
  wire [63:0] _895;
  wire [63:0] _894;
  wire [63:0] _893;
  wire [63:0] _892;
  wire [63:0] _891;
  wire [63:0] _890;
  wire [63:0] _889;
  wire [63:0] _888;
  wire [63:0] _887;
  wire [63:0] _886;
  wire [63:0] _885;
  wire [63:0] _884;
  wire [63:0] _883;
  wire [63:0] _882;
  wire [63:0] _881;
  wire [63:0] _880;
  wire [63:0] _879;
  wire [63:0] _878;
  wire [63:0] _877;
  wire [31:0] _876;
  wire [63:0] _875;
  wire [63:0] _874;
  wire [63:0] _873;
  wire [0:0] ifout903;
  wire [63:0] _872;
  wire [63:0] _871;
  wire [63:0] _870;
  wire [63:0] _869;
  wire [63:0] _868;
  wire [63:0] _867;
  wire [31:0] off_3611;
  wire [31:0] _866;
  wire [63:0] _865;
  wire [31:0] idx_3610;
  wire [31:0] _864;
  wire [31:0] _863;
  wire [63:0] _862;
  wire [63:0] _861;
  wire [63:0] _860;
  wire [63:0] _859;
  wire [63:0] _858;
  wire [63:0] _857;
  wire [63:0] _856;
  wire [63:0] _855;
  wire [63:0] _854;
  wire [63:0] _853;
  wire [63:0] _852;
  wire [63:0] _851;
  wire [63:0] _850;
  wire [63:0] _849;
  wire [63:0] _848;
  wire [63:0] _847;
  wire [63:0] _846;
  wire [63:0] _845;
  wire [63:0] _844;
  wire [63:0] _843;
  wire [63:0] _842;
  wire [63:0] _841;
  wire [63:0] _840;
  wire [63:0] _839;
  wire [63:0] _838;
  wire [63:0] _837;
  wire [63:0] _836;
  wire [63:0] _835;
  wire [63:0] _834;
  wire [63:0] _833;
  wire [63:0] _832;
  wire [63:0] _831;
  wire [63:0] _830;
  wire [63:0] _829;
  wire [63:0] _828;
  wire [63:0] _827;
  wire [63:0] _826;
  wire [63:0] _825;
  wire [63:0] _824;
  wire [63:0] _823;
  wire [63:0] _822;
  wire [63:0] _821;
  wire [63:0] _820;
  wire [63:0] _819;
  wire [63:0] _818;
  wire [63:0] _817;
  wire [63:0] _816;
  wire [63:0] _815;
  wire [63:0] _814;
  wire [63:0] _813;
  wire [63:0] _812;
  wire [63:0] _811;
  wire [63:0] _810;
  wire [63:0] _809;
  wire [63:0] _808;
  wire [63:0] _807;
  wire [63:0] _806;
  wire [63:0] _805;
  wire [63:0] _804;
  wire [63:0] _803;
  wire [63:0] _802;
  wire [63:0] _801;
  wire [63:0] _800;
  wire [63:0] _799;
  wire [63:0] _798;
  wire [63:0] _797;
  wire [63:0] _796;
  wire [63:0] _795;
  wire [63:0] _794;
  wire [63:0] _793;
  wire [63:0] _792;
  wire [63:0] _791;
  wire [63:0] _790;
  wire [63:0] _789;
  wire [63:0] _788;
  wire [63:0] _787;
  wire [63:0] _786;
  wire [63:0] _785;
  wire [63:0] _784;
  wire [63:0] _783;
  wire [63:0] _782;
  wire [31:0] _781;
  wire [63:0] _780;
  wire [63:0] _779;
  wire [63:0] _778;
  wire [0:0] ifout805;
  wire [63:0] _777;
  wire [63:0] _776;
  wire [63:0] _775;
  wire [63:0] _774;
  wire [63:0] _773;
  wire [63:0] _772;
  wire [31:0] off_3603;
  wire [63:0] _771;
  wire [31:0] idx_3601;
  wire [31:0] _770;
  wire [31:0] _769;
  wire [63:0] _768;
  wire [63:0] _767;
  wire [63:0] _766;
  wire [63:0] _765;
  wire [63:0] _764;
  wire [63:0] _763;
  wire [63:0] _762;
  wire [63:0] _761;
  wire [63:0] _760;
  wire [63:0] _759;
  wire [63:0] _758;
  wire [63:0] _757;
  wire [63:0] _756;
  wire [63:0] _755;
  wire [63:0] _754;
  wire [63:0] _753;
  wire [63:0] _752;
  wire [63:0] _751;
  wire [63:0] _750;
  wire [63:0] _749;
  wire [63:0] _748;
  wire [63:0] _747;
  wire [63:0] _746;
  wire [63:0] _745;
  wire [63:0] _744;
  wire [63:0] _743;
  wire [63:0] _742;
  wire [63:0] _741;
  wire [63:0] _740;
  wire [63:0] _739;
  wire [63:0] _738;
  wire [63:0] _737;
  wire [63:0] _736;
  wire [63:0] _735;
  wire [63:0] _734;
  wire [63:0] _733;
  wire [63:0] _732;
  wire [63:0] _731;
  wire [63:0] _730;
  wire [63:0] _729;
  wire [63:0] _728;
  wire [63:0] _727;
  wire [63:0] _726;
  wire [63:0] _725;
  wire [63:0] _724;
  wire [63:0] _723;
  wire [63:0] _722;
  wire [63:0] _721;
  wire [63:0] _720;
  wire [63:0] _719;
  wire [63:0] _718;
  wire [63:0] _717;
  wire [63:0] _716;
  wire [63:0] _715;
  wire [63:0] _714;
  wire [63:0] _713;
  wire [63:0] _712;
  wire [63:0] _711;
  wire [63:0] _710;
  wire [63:0] _709;
  wire [63:0] _708;
  wire [63:0] _707;
  wire [63:0] _706;
  wire [63:0] _705;
  wire [63:0] _704;
  wire [63:0] _703;
  wire [63:0] _702;
  wire [63:0] _701;
  wire [63:0] _700;
  wire [63:0] _699;
  wire [63:0] _698;
  wire [63:0] _697;
  wire [63:0] _696;
  wire [63:0] _695;
  wire [63:0] _694;
  wire [63:0] _693;
  wire [63:0] _692;
  wire [63:0] _691;
  wire [63:0] _690;
  wire [63:0] _689;
  wire [63:0] _688;
  wire [31:0] _687;
  wire [63:0] _686;
  wire [63:0] _685;
  wire [63:0] _684;
  wire [0:0] ifout708;
  wire [63:0] _683;
  wire [63:0] _682;
  wire [63:0] _681;
  wire [63:0] _680;
  wire [63:0] _679;
  wire [63:0] _678;
  wire [31:0] off_3594;
  wire [31:0] _677;
  wire [31:0] idx_3593;
  wire [31:0] _676;
  wire [31:0] _675;
  wire [63:0] _674;
  wire [63:0] _673;
  wire [63:0] _672;
  wire [63:0] _671;
  wire [63:0] _670;
  wire [63:0] _669;
  wire [63:0] _668;
  wire [63:0] _667;
  wire [63:0] _666;
  wire [63:0] _665;
  wire [63:0] _664;
  wire [63:0] _663;
  wire [63:0] _662;
  wire [63:0] _661;
  wire [63:0] _660;
  wire [63:0] _659;
  wire [63:0] _658;
  wire [63:0] _657;
  wire [63:0] _656;
  wire [63:0] _655;
  wire [63:0] _654;
  wire [63:0] _653;
  wire [63:0] _652;
  wire [63:0] _651;
  wire [63:0] _650;
  wire [63:0] _649;
  wire [63:0] _648;
  wire [63:0] _647;
  wire [63:0] _646;
  wire [63:0] _645;
  wire [63:0] _644;
  wire [63:0] _643;
  wire [63:0] _642;
  wire [63:0] _641;
  wire [63:0] _640;
  wire [63:0] _639;
  wire [63:0] _638;
  wire [63:0] _637;
  wire [63:0] _636;
  wire [63:0] _635;
  wire [63:0] _634;
  wire [63:0] _633;
  wire [63:0] _632;
  wire [63:0] _631;
  wire [63:0] _630;
  wire [63:0] _629;
  wire [63:0] _628;
  wire [63:0] _627;
  wire [63:0] _626;
  wire [63:0] _625;
  wire [63:0] _624;
  wire [63:0] _623;
  wire [63:0] _622;
  wire [63:0] _621;
  wire [63:0] _620;
  wire [63:0] _619;
  wire [63:0] _618;
  wire [63:0] _617;
  wire [63:0] _616;
  wire [63:0] _615;
  wire [63:0] _614;
  wire [63:0] _613;
  wire [63:0] _612;
  wire [63:0] _611;
  wire [63:0] _610;
  wire [63:0] _609;
  wire [63:0] _608;
  wire [63:0] _607;
  wire [63:0] _606;
  wire [63:0] _605;
  wire [63:0] _604;
  wire [63:0] _603;
  wire [63:0] _602;
  wire [63:0] _601;
  wire [63:0] _600;
  wire [63:0] _599;
  wire [63:0] _598;
  wire [63:0] _597;
  wire [63:0] _596;
  wire [63:0] _595;
  wire [63:0] _594;
  wire [31:0] _593;
  wire [63:0] _592;
  wire [63:0] _591;
  wire [63:0] _590;
  wire [0:0] ifout611;
  wire [63:0] _589;
  wire [63:0] _588;
  wire [63:0] _587;
  wire [63:0] _586;
  wire [63:0] _585;
  wire [63:0] _584;
  wire [31:0] off_3586;
  wire [31:0] _583;
  wire [63:0] _582;
  wire [31:0] idx_3585;
  wire [31:0] _581;
  wire [31:0] _580;
  wire [63:0] _579;
  wire [63:0] _578;
  wire [63:0] _577;
  wire [63:0] _576;
  wire [63:0] _575;
  wire [63:0] _574;
  wire [63:0] _573;
  wire [63:0] _572;
  wire [63:0] _571;
  wire [63:0] _570;
  wire [63:0] _569;
  wire [63:0] _568;
  wire [63:0] _567;
  wire [63:0] _566;
  wire [63:0] _565;
  wire [63:0] _564;
  wire [63:0] _563;
  wire [63:0] _562;
  wire [63:0] _561;
  wire [63:0] _560;
  wire [63:0] _559;
  wire [63:0] _558;
  wire [63:0] _557;
  wire [63:0] _556;
  wire [63:0] _555;
  wire [63:0] _554;
  wire [63:0] _553;
  wire [63:0] _552;
  wire [63:0] _551;
  wire [63:0] _550;
  wire [63:0] _549;
  wire [63:0] _548;
  wire [63:0] _547;
  wire [63:0] _546;
  wire [63:0] _545;
  wire [63:0] _544;
  wire [63:0] _543;
  wire [63:0] _542;
  wire [63:0] _541;
  wire [63:0] _540;
  wire [63:0] _539;
  wire [63:0] _538;
  wire [63:0] _537;
  wire [63:0] _536;
  wire [63:0] _535;
  wire [63:0] _534;
  wire [63:0] _533;
  wire [63:0] _532;
  wire [63:0] _531;
  wire [63:0] _530;
  wire [63:0] _529;
  wire [63:0] _528;
  wire [63:0] _527;
  wire [63:0] _526;
  wire [63:0] _525;
  wire [63:0] _524;
  wire [63:0] _523;
  wire [63:0] _522;
  wire [63:0] _521;
  wire [63:0] _520;
  wire [63:0] _519;
  wire [63:0] _518;
  wire [63:0] _517;
  wire [63:0] _516;
  wire [63:0] _515;
  wire [63:0] _514;
  wire [63:0] _513;
  wire [63:0] _512;
  wire [63:0] _511;
  wire [63:0] _510;
  wire [63:0] _509;
  wire [63:0] _508;
  wire [63:0] _507;
  wire [63:0] _506;
  wire [63:0] _505;
  wire [63:0] _504;
  wire [63:0] _503;
  wire [63:0] _502;
  wire [63:0] _501;
  wire [63:0] _500;
  wire [63:0] _499;
  wire [31:0] _498;
  wire [63:0] _497;
  wire [63:0] _496;
  wire [63:0] _495;
  wire [0:0] ifout513;
  wire [63:0] _494;
  wire [63:0] _493;
  wire [63:0] _492;
  wire [63:0] _491;
  wire [63:0] _490;
  wire [63:0] _489;
  wire [31:0] off_3578;
  wire [31:0] _488;
  wire [63:0] _487;
  wire [31:0] idx_3577;
  wire [31:0] _486;
  wire [31:0] _485;
  wire [63:0] _484;
  wire [63:0] _483;
  wire [63:0] _482;
  wire [63:0] _481;
  wire [63:0] _480;
  wire [63:0] _479;
  wire [63:0] _478;
  wire [63:0] _477;
  wire [63:0] _476;
  wire [63:0] _475;
  wire [63:0] _474;
  wire [63:0] _473;
  wire [63:0] _472;
  wire [63:0] _471;
  wire [63:0] _470;
  wire [63:0] _469;
  wire [63:0] _468;
  wire [63:0] _467;
  wire [63:0] _466;
  wire [63:0] _465;
  wire [63:0] _464;
  wire [63:0] _463;
  wire [63:0] _462;
  wire [63:0] _461;
  wire [63:0] _460;
  wire [63:0] _459;
  wire [63:0] _458;
  wire [63:0] _457;
  wire [63:0] _456;
  wire [63:0] _455;
  wire [63:0] _454;
  wire [63:0] _453;
  wire [63:0] _452;
  wire [63:0] _451;
  wire [63:0] _450;
  wire [63:0] _449;
  wire [63:0] _448;
  wire [63:0] _447;
  wire [63:0] _446;
  wire [63:0] _445;
  wire [63:0] _444;
  wire [63:0] _443;
  wire [63:0] _442;
  wire [63:0] _441;
  wire [63:0] _440;
  wire [63:0] _439;
  wire [63:0] _438;
  wire [63:0] _437;
  wire [63:0] _436;
  wire [63:0] _435;
  wire [63:0] _434;
  wire [63:0] _433;
  wire [63:0] _432;
  wire [63:0] _431;
  wire [63:0] _430;
  wire [63:0] _429;
  wire [63:0] _428;
  wire [63:0] _427;
  wire [63:0] _426;
  wire [63:0] _425;
  wire [63:0] _424;
  wire [63:0] _423;
  wire [63:0] _422;
  wire [63:0] _421;
  wire [63:0] _420;
  wire [63:0] _419;
  wire [63:0] _418;
  wire [63:0] _417;
  wire [63:0] _416;
  wire [63:0] _415;
  wire [63:0] _414;
  wire [63:0] _413;
  wire [63:0] _412;
  wire [63:0] _411;
  wire [63:0] _410;
  wire [63:0] _409;
  wire [63:0] _408;
  wire [63:0] _407;
  wire [63:0] _406;
  wire [63:0] _405;
  wire [63:0] _404;
  wire [31:0] _403;
  wire [63:0] _402;
  wire [63:0] _401;
  wire [63:0] _400;
  wire [0:0] ifout415;
  wire [63:0] _399;
  wire [63:0] _398;
  wire [63:0] _397;
  wire [63:0] _396;
  wire [63:0] _395;
  wire [63:0] _394;
  wire [31:0] off_3570;
  wire [31:0] _393;
  wire [63:0] _392;
  wire [31:0] idx_3569;
  wire [31:0] _391;
  wire [31:0] _390;
  wire [63:0] _389;
  wire [63:0] _388;
  wire [63:0] _387;
  wire [63:0] _386;
  wire [63:0] _385;
  wire [63:0] _384;
  wire [63:0] _383;
  wire [63:0] _382;
  wire [63:0] _381;
  wire [63:0] _380;
  wire [63:0] _379;
  wire [63:0] _378;
  wire [63:0] _377;
  wire [63:0] _376;
  wire [63:0] _375;
  wire [63:0] _374;
  wire [63:0] _373;
  wire [63:0] _372;
  wire [63:0] _371;
  wire [63:0] _370;
  wire [63:0] _369;
  wire [63:0] _368;
  wire [63:0] _367;
  wire [63:0] _366;
  wire [63:0] _365;
  wire [63:0] _364;
  wire [63:0] _363;
  wire [63:0] _362;
  wire [63:0] _361;
  wire [63:0] _360;
  wire [63:0] _359;
  wire [63:0] _358;
  wire [63:0] _357;
  wire [63:0] _356;
  wire [63:0] _355;
  wire [63:0] _354;
  wire [63:0] _353;
  wire [63:0] _352;
  wire [63:0] _351;
  wire [63:0] _350;
  wire [63:0] _349;
  wire [63:0] _348;
  wire [63:0] _347;
  wire [63:0] _346;
  wire [63:0] _345;
  wire [63:0] _344;
  wire [63:0] _343;
  wire [63:0] _342;
  wire [63:0] _341;
  wire [63:0] _340;
  wire [63:0] _339;
  wire [63:0] _338;
  wire [63:0] _337;
  wire [63:0] _336;
  wire [63:0] _335;
  wire [63:0] _334;
  wire [63:0] _333;
  wire [63:0] _332;
  wire [63:0] _331;
  wire [63:0] _330;
  wire [63:0] _329;
  wire [63:0] _328;
  wire [63:0] _327;
  wire [63:0] _326;
  wire [63:0] _325;
  wire [63:0] _324;
  wire [63:0] _323;
  wire [63:0] _322;
  wire [63:0] _321;
  wire [63:0] _320;
  wire [63:0] _319;
  wire [63:0] _318;
  wire [63:0] _317;
  wire [63:0] _316;
  wire [63:0] _315;
  wire [63:0] _314;
  wire [63:0] _313;
  wire [63:0] _312;
  wire [63:0] _311;
  wire [63:0] _310;
  wire [63:0] _309;
  wire [31:0] _308;
  wire [63:0] _307;
  wire [63:0] _306;
  wire [63:0] _305;
  wire [0:0] ifout317;
  wire [63:0] _304;
  wire [63:0] _303;
  wire [63:0] _302;
  wire [63:0] _301;
  wire [63:0] _300;
  wire [63:0] _299;
  wire [31:0] off_3562;
  wire [31:0] _298;
  wire [63:0] _297;
  wire [31:0] idx_3561;
  wire [31:0] _296;
  wire [31:0] _295;
  wire [63:0] _294;
  wire [63:0] _293;
  wire [63:0] _292;
  wire [63:0] _291;
  wire [63:0] _290;
  wire [63:0] _289;
  wire [63:0] _288;
  wire [63:0] _287;
  wire [63:0] _286;
  wire [63:0] _285;
  wire [63:0] _284;
  wire [63:0] _283;
  wire [63:0] _282;
  wire [63:0] _281;
  wire [63:0] _280;
  wire [63:0] _279;
  wire [63:0] _278;
  wire [63:0] _277;
  wire [63:0] _276;
  wire [63:0] _275;
  wire [63:0] _274;
  wire [63:0] _273;
  wire [63:0] _272;
  wire [63:0] _271;
  wire [63:0] _270;
  wire [63:0] _269;
  wire [63:0] _268;
  wire [63:0] _267;
  wire [63:0] _266;
  wire [63:0] _265;
  wire [63:0] _264;
  wire [63:0] _263;
  wire [63:0] _262;
  wire [63:0] _261;
  wire [63:0] _260;
  wire [63:0] _259;
  wire [63:0] _258;
  wire [63:0] _257;
  wire [63:0] _256;
  wire [63:0] _255;
  wire [63:0] _254;
  wire [63:0] _253;
  wire [63:0] _252;
  wire [63:0] _251;
  wire [63:0] _250;
  wire [63:0] _249;
  wire [63:0] _248;
  wire [63:0] _247;
  wire [63:0] _246;
  wire [63:0] _245;
  wire [63:0] _244;
  wire [63:0] _243;
  wire [63:0] _242;
  wire [63:0] _241;
  wire [63:0] _240;
  wire [63:0] _239;
  wire [63:0] _238;
  wire [63:0] _237;
  wire [63:0] _236;
  wire [63:0] _235;
  wire [63:0] _234;
  wire [63:0] _233;
  wire [63:0] _232;
  wire [63:0] _231;
  wire [63:0] _230;
  wire [63:0] _229;
  wire [63:0] _228;
  wire [63:0] _227;
  wire [63:0] _226;
  wire [63:0] _225;
  wire [63:0] _224;
  wire [63:0] _223;
  wire [63:0] _222;
  wire [63:0] _221;
  wire [63:0] _220;
  wire [63:0] _219;
  wire [63:0] _218;
  wire [63:0] _217;
  wire [63:0] _216;
  wire [63:0] _215;
  wire [63:0] _214;
  wire [31:0] _213;
  wire [63:0] _212;
  wire [63:0] _211;
  wire [63:0] _210;
  wire [0:0] ifout219;
  wire [63:0] _209;
  wire [63:0] _208;
  wire [63:0] _207;
  wire [63:0] _206;
  wire [63:0] _205;
  wire [63:0] _204;
  wire [31:0] off_3554;
  wire [31:0] _203;
  wire [63:0] _202;
  wire [31:0] idx_3553;
  wire [31:0] _201;
  wire [31:0] _200;
  wire [63:0] _199;
  wire [63:0] _198;
  wire [63:0] _197;
  wire [63:0] _196;
  wire [63:0] _195;
  wire [63:0] _194;
  wire [63:0] _193;
  wire [63:0] _192;
  wire [63:0] _191;
  wire [63:0] _190;
  wire [63:0] _189;
  wire [63:0] _188;
  wire [63:0] _187;
  wire [63:0] _186;
  wire [63:0] _185;
  wire [63:0] _184;
  wire [63:0] _183;
  wire [63:0] _182;
  wire [63:0] _181;
  wire [63:0] _180;
  wire [63:0] _179;
  wire [63:0] _178;
  wire [63:0] _177;
  wire [63:0] _176;
  wire [63:0] _175;
  wire [63:0] _174;
  wire [63:0] _173;
  wire [63:0] _172;
  wire [63:0] _171;
  wire [63:0] _170;
  wire [63:0] _169;
  wire [63:0] _168;
  wire [63:0] _167;
  wire [63:0] _166;
  wire [63:0] _165;
  wire [63:0] _164;
  wire [63:0] _163;
  wire [63:0] _162;
  wire [63:0] _161;
  wire [63:0] _160;
  wire [63:0] _159;
  wire [63:0] _158;
  wire [63:0] _157;
  wire [63:0] _156;
  wire [63:0] _155;
  wire [63:0] _154;
  wire [63:0] _153;
  wire [63:0] _152;
  wire [63:0] _151;
  wire [63:0] _150;
  wire [63:0] _149;
  wire [63:0] _148;
  wire [63:0] _147;
  wire [63:0] _146;
  wire [63:0] _145;
  wire [63:0] _144;
  wire [63:0] _143;
  wire [63:0] _142;
  wire [63:0] _141;
  wire [63:0] _140;
  wire [63:0] _139;
  wire [63:0] _138;
  wire [63:0] _137;
  wire [63:0] _136;
  wire [63:0] _135;
  wire [63:0] _134;
  wire [63:0] _133;
  wire [63:0] _132;
  wire [63:0] _131;
  wire [63:0] _130;
  wire [63:0] _129;
  wire [63:0] _128;
  wire [63:0] _127;
  wire [63:0] _126;
  wire [63:0] _125;
  wire [63:0] _124;
  wire [63:0] _123;
  wire [63:0] _122;
  wire [63:0] _121;
  wire [63:0] _120;
  wire [63:0] _119;
  wire [31:0] _118;
  wire [63:0] _117;
  wire [63:0] _116;
  wire [63:0] _115;
  wire [0:0] ifout121;
  wire [63:0] _114;
  wire [63:0] _113;
  wire [63:0] _112;
  wire [63:0] _111;
  wire [63:0] _110;
  wire [63:0] _109;
  wire [31:0] off_3546;
  wire [31:0] _108;
  wire [63:0] _107;
  wire [31:0] idx_3545;
  wire [31:0] _106;
  wire [31:0] _105;
  wire [63:0] _104;
  wire [63:0] _103;
  wire [63:0] _102;
  wire [63:0] _101;
  wire [63:0] _100;
  wire [63:0] _99;
  wire [63:0] _98;
  wire [63:0] _97;
  wire [63:0] _96;
  wire [63:0] _95;
  wire [63:0] _94;
  wire [63:0] _93;
  wire [63:0] _92;
  wire [63:0] _91;
  wire [63:0] _90;
  wire [63:0] _89;
  wire [63:0] _88;
  wire [63:0] _87;
  wire [63:0] _86;
  wire [63:0] _85;
  wire [63:0] _84;
  wire [63:0] _83;
  wire [63:0] _82;
  wire [63:0] _81;
  wire [63:0] _80;
  wire [63:0] _79;
  wire [63:0] _78;
  wire [63:0] _77;
  wire [63:0] _76;
  wire [63:0] _75;
  wire [63:0] _74;
  wire [63:0] _73;
  wire [63:0] _72;
  wire [63:0] _71;
  wire [63:0] _70;
  wire [63:0] _69;
  wire [63:0] _68;
  wire [63:0] _67;
  wire [63:0] _66;
  wire [63:0] _65;
  wire [63:0] _64;
  wire [63:0] _63;
  wire [63:0] _62;
  wire [63:0] _61;
  wire [63:0] _60;
  wire [63:0] _59;
  wire [63:0] _58;
  wire [63:0] _57;
  wire [63:0] _56;
  wire [63:0] _55;
  wire [63:0] _54;
  wire [63:0] _53;
  wire [63:0] _52;
  wire [63:0] _51;
  wire [63:0] _50;
  wire [63:0] _49;
  wire [63:0] _48;
  wire [63:0] _47;
  wire [63:0] _46;
  wire [63:0] _45;
  wire [63:0] _44;
  wire [63:0] _43;
  wire [63:0] _42;
  wire [63:0] _41;
  wire [63:0] _40;
  wire [63:0] _39;
  wire [63:0] _38;
  wire [63:0] _37;
  wire [63:0] _36;
  wire [63:0] _35;
  wire [63:0] _34;
  wire [63:0] _33;
  wire [63:0] _32;
  wire [63:0] _31;
  wire [63:0] _30;
  wire [63:0] _29;
  wire [63:0] _28;
  wire [63:0] _27;
  wire [63:0] _26;
  wire [63:0] _25;
  wire [63:0] _24;
  wire [31:0] _23;
  wire [63:0] _22;
  wire [63:0] _21;
  wire [63:0] _20;
  wire [0:0] ifout23;
  wire [63:0] _19;
  wire [63:0] _18;
  wire [63:0] _17;
  wire [63:0] _16;
  wire [63:0] _15;
  wire [63:0] _14;
  wire [31:0] off_3537;
  wire [31:0] _13;
  wire [63:0] _12;
  wire [31:0] idx_3536;
  wire [31:0] _11;
  wire [31:0] _10;
  wire [15:0] _9;
  wire [63:0] _8;
  wire [63:0] _7;
  wire [63:0] _6;
  wire [0:0] ifout6;
  wire [15:0] _5;
  wire [63:0] _4;
  wire [63:0] _3;
  wire [63:0] _2;
  wire [31:0] idx_3531;
  wire [63:0] _1;
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op0 (.out1(_1), .in1(ip1_3530_D), .in2(6 'd 48));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1 (.out1(idx_3531), .in1(_1));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3683 (.out1(R3684), .clock(clock), .in1(idx_3531));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2 (.out1(_2), .in1(R3684));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op3 (.out1(_3), .in1(_2), .in2(1 'd 1));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3684 (.out1(R3685), .clock(clock), .in1(R3684));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3940 (.out1(R3941), .clock(clock), .in1(_3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op4 (.out1(_4), .in1(dirC_3532_D), .in2(R3941));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3685 (.out1(R3686), .clock(clock), .in1(R3685));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op3941 (.out1(R3942), .clock(clock), .in1(_4));
  SRAM op5 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_5),.ADR(R3942));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3686 (.out1(R3687), .clock(clock), .in1(R3686));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op3942 (.out1(R3943), .clock(clock), .in1(_5));
  NE_EXPR #(.BITSIZE_in1(16), .BITSIZE_in2(1),.BITSIZE_out1(1)) op6 (.out1(ifout6), .in1(R3943), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op7 (.out1(_6), .in1(R3687));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op8 (.out1(_7), .in1(_6), .in2(1 'd 1));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3687 (.out1(R3688), .clock(clock), .in1(R3687));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3943 (.out1(R3944), .clock(clock), .in1(ifout6));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4198 (.out1(R4199), .clock(clock), .in1(_7));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op9 (.out1(_8), .in1(dirC_3532_D), .in2(R4199));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3688 (.out1(R3689), .clock(clock), .in1(R3688));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3944 (.out1(R3945), .clock(clock), .in1(R3944));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4199 (.out1(R4200), .clock(clock), .in1(_8));
  SRAM op10 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_9),.ADR(R4200));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3689 (.out1(R3690), .clock(clock), .in1(R3689));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3945 (.out1(R3946), .clock(clock), .in1(R3945));
  REG_STD #(.BITSIZE_in1(16), .BITSIZE_out1(16)) op4200 (.out1(R4201), .clock(clock), .in1(_9));
  cast #(.BITSIZE_in1(16), .BITSIZE_out1(32)) op11 (.out1(_10), .in1(R4201));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(1), .BITSIZE_out1(32)) op12 (.out1(_11), .in1(_10), .in2(-1 'd 1));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13 (.out1(idx_3536), .in1(_11));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3690 (.out1(R3691), .clock(clock), .in1(R3690));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3946 (.out1(R3947), .clock(clock), .in1(R3946));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4201 (.out1(R4202), .clock(clock), .in1(idx_3536));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op17 (.out1(_14), .in1(R4202));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op18 (.out1(_15), .in1(_14), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3691 (.out1(R3692), .clock(clock), .in1(R3691));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3947 (.out1(R3948), .clock(clock), .in1(R3947));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4202 (.out1(R4203), .clock(clock), .in1(R4202));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4447 (.out1(R4448), .clock(clock), .in1(_15));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op19 (.out1(_16), .in1(vec16_3538_D), .in2(R4448));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3692 (.out1(R3693), .clock(clock), .in1(R3692));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3948 (.out1(R3949), .clock(clock), .in1(R3948));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4203 (.out1(R4204), .clock(clock), .in1(R4203));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4448 (.out1(R4449), .clock(clock), .in1(_16));
  SRAM op20 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_17),.ADR(R4449));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3693 (.out1(R3694), .clock(clock), .in1(R3693));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3949 (.out1(R3950), .clock(clock), .in1(R3949));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4204 (.out1(R4205), .clock(clock), .in1(R4204));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4449 (.out1(R4450), .clock(clock), .in1(_17));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op14 (.out1(_12), .in1(ip1_3530_D), .in2(6 'd 42));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op15 (.out1(_13), .in1(_12));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op16 (.out1(off_3537), .in1(_13), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op21 (.out1(_18), .in1(R4450), .in2(off_3537));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3694 (.out1(R3695), .clock(clock), .in1(R3694));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3950 (.out1(R3951), .clock(clock), .in1(R3950));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4205 (.out1(R4206), .clock(clock), .in1(R4205));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4450 (.out1(R4451), .clock(clock), .in1(off_3537));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4690 (.out1(R4691), .clock(clock), .in1(_18));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op22 (.out1(_19), .in1(R4691), .in2(1 'd 1));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op23 (.out1(ifout23), .in1(_19), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op91 (.out1(_87), .in1(R4206));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op84 (.out1(_80), .in1(R4206));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op73 (.out1(_69), .in1(R4206));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op53 (.out1(_49), .in1(R4206));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op92 (.out1(_88), .in1(_87), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op85 (.out1(_81), .in1(_80), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op74 (.out1(_70), .in1(_69), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op54 (.out1(_50), .in1(_49), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3695 (.out1(R3696), .clock(clock), .in1(R3695));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3951 (.out1(R3952), .clock(clock), .in1(R3951));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4206 (.out1(R4207), .clock(clock), .in1(R4206));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4451 (.out1(R4452), .clock(clock), .in1(R4451));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4691 (.out1(R4692), .clock(clock), .in1(ifout23));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4938 (.out1(R4939), .clock(clock), .in1(_88));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4939 (.out1(R4940), .clock(clock), .in1(_81));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4940 (.out1(R4941), .clock(clock), .in1(_70));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4941 (.out1(R4942), .clock(clock), .in1(_50));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op66 (.out1(_62), .in1(R4207));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op46 (.out1(_42), .in1(R4207));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op35 (.out1(_31), .in1(R4207));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op28 (.out1(_24), .in1(R4207));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op95 (.out1(_91), .in1(2 'd 2), .in2(R4452));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op67 (.out1(_63), .in1(_62), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op47 (.out1(_43), .in1(_42), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op36 (.out1(_32), .in1(_31), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op29 (.out1(_25), .in1(_24), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op93 (.out1(_89), .in1(vec16_3538_D), .in2(R4939));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op86 (.out1(_82), .in1(vec16_3538_D), .in2(R4940));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op75 (.out1(_71), .in1(vec16_3538_D), .in2(R4941));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op55 (.out1(_51), .in1(vec16_3538_D), .in2(R4942));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3696 (.out1(R3697), .clock(clock), .in1(R3696));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3952 (.out1(R3953), .clock(clock), .in1(R3952));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4207 (.out1(R4208), .clock(clock), .in1(R4207));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4452 (.out1(R4453), .clock(clock), .in1(R4452));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4692 (.out1(R4693), .clock(clock), .in1(R4692));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4942 (.out1(R4943), .clock(clock), .in1(_91));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4943 (.out1(R4944), .clock(clock), .in1(_63));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4944 (.out1(R4945), .clock(clock), .in1(_43));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4945 (.out1(R4946), .clock(clock), .in1(_32));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4946 (.out1(R4947), .clock(clock), .in1(_25));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4947 (.out1(R4948), .clock(clock), .in1(_89));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4948 (.out1(R4949), .clock(clock), .in1(_82));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4949 (.out1(R4950), .clock(clock), .in1(_71));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4950 (.out1(R4951), .clock(clock), .in1(_51));
  SRAM op94 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_90),.ADR(R4948));
  SRAM op87 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_83),.ADR(R4949));
  SRAM op76 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_72),.ADR(R4950));
  SRAM op56 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_52),.ADR(R4951));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op88 (.out1(_84), .in1(2 'd 2), .in2(R4453));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op77 (.out1(_73), .in1(2 'd 2), .in2(R4453));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op70 (.out1(_66), .in1(2 'd 2), .in2(R4453));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op57 (.out1(_53), .in1(2 'd 2), .in2(R4453));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op50 (.out1(_46), .in1(2 'd 2), .in2(R4453));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op39 (.out1(_35), .in1(2 'd 2), .in2(R4453));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op68 (.out1(_64), .in1(vec16_3538_D), .in2(R4944));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op48 (.out1(_44), .in1(vec16_3538_D), .in2(R4945));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op37 (.out1(_33), .in1(vec16_3538_D), .in2(R4946));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op30 (.out1(_26), .in1(vec16_3538_D), .in2(R4947));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op96 (.out1(_92), .in1(R4943), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3697 (.out1(R3698), .clock(clock), .in1(R3697));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3953 (.out1(R3954), .clock(clock), .in1(R3953));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4208 (.out1(R4209), .clock(clock), .in1(R4208));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4453 (.out1(R4454), .clock(clock), .in1(R4453));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4693 (.out1(R4694), .clock(clock), .in1(R4693));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4951 (.out1(R4952), .clock(clock), .in1(_90));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4952 (.out1(R4953), .clock(clock), .in1(_83));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4953 (.out1(R4954), .clock(clock), .in1(_72));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4954 (.out1(R4955), .clock(clock), .in1(_52));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4955 (.out1(R4956), .clock(clock), .in1(_84));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4956 (.out1(R4957), .clock(clock), .in1(_73));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4957 (.out1(R4958), .clock(clock), .in1(_66));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4958 (.out1(R4959), .clock(clock), .in1(_53));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4959 (.out1(R4960), .clock(clock), .in1(_46));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4960 (.out1(R4961), .clock(clock), .in1(_35));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4961 (.out1(R4962), .clock(clock), .in1(_64));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4962 (.out1(R4963), .clock(clock), .in1(_44));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4963 (.out1(R4964), .clock(clock), .in1(_33));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4964 (.out1(R4965), .clock(clock), .in1(_26));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4965 (.out1(R4966), .clock(clock), .in1(_92));
  SRAM op69 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_65),.ADR(R4962));
  SRAM op49 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_45),.ADR(R4963));
  SRAM op38 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_34),.ADR(R4964));
  SRAM op31 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_27),.ADR(R4965));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op97 (.out1(_93), .in1(R4952), .in2(R4966));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op98 (.out1(_94), .in1(_93), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op89 (.out1(_85), .in1(R4956), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op78 (.out1(_74), .in1(R4957), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op58 (.out1(_54), .in1(R4959), .in2(64 'd 18446744073709551615));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op32 (.out1(_28), .in1(2 'd 2), .in2(R4454));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op99 (.out1(_95), .in1(_94), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op90 (.out1(_86), .in1(R4953), .in2(_85));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op79 (.out1(_75), .in1(R4954), .in2(_74));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op59 (.out1(_55), .in1(R4955), .in2(_54));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op100 (.out1(_96), .in1(_86), .in2(_95));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op80 (.out1(_76), .in1(_75), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op71 (.out1(_67), .in1(R4958), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op60 (.out1(_56), .in1(_55), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op51 (.out1(_47), .in1(R4960), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op40 (.out1(_36), .in1(R4961), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3698 (.out1(R3699), .clock(clock), .in1(R3698));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3954 (.out1(R3955), .clock(clock), .in1(R3954));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4209 (.out1(R4210), .clock(clock), .in1(R4209));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4454 (.out1(R4455), .clock(clock), .in1(R4454));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4694 (.out1(R4695), .clock(clock), .in1(R4694));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4966 (.out1(R4967), .clock(clock), .in1(_65));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4967 (.out1(R4968), .clock(clock), .in1(_45));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4968 (.out1(R4969), .clock(clock), .in1(_34));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4969 (.out1(R4970), .clock(clock), .in1(_27));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4970 (.out1(R4971), .clock(clock), .in1(_28));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4971 (.out1(R4972), .clock(clock), .in1(_96));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4972 (.out1(R4973), .clock(clock), .in1(_76));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4973 (.out1(R4974), .clock(clock), .in1(_67));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4974 (.out1(R4975), .clock(clock), .in1(_56));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4975 (.out1(R4976), .clock(clock), .in1(_47));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4976 (.out1(R4977), .clock(clock), .in1(_36));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op81 (.out1(_77), .in1(R4973), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op72 (.out1(_68), .in1(R4967), .in2(R4974));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op41 (.out1(_37), .in1(R4969), .in2(R4977));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op101 (.out1(_97), .in1(R4972), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op82 (.out1(_78), .in1(_68), .in2(_77));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op61 (.out1(_57), .in1(R4975), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op52 (.out1(_48), .in1(R4968), .in2(R4976));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op42 (.out1(_38), .in1(_37), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op33 (.out1(_29), .in1(R4971), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op62 (.out1(_58), .in1(_48), .in2(_57));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op102 (.out1(_98), .in1(_97), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op83 (.out1(_79), .in1(_78), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op43 (.out1(_39), .in1(_38), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op34 (.out1(_30), .in1(R4970), .in2(_29));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op103 (.out1(_99), .in1(_79), .in2(_98));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op63 (.out1(_59), .in1(_58), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op44 (.out1(_40), .in1(_30), .in2(_39));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3699 (.out1(R3700), .clock(clock), .in1(R3699));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3955 (.out1(R3956), .clock(clock), .in1(R3955));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4210 (.out1(R4211), .clock(clock), .in1(R4210));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4455 (.out1(R4456), .clock(clock), .in1(R4455));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4695 (.out1(R4696), .clock(clock), .in1(R4695));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4977 (.out1(R4978), .clock(clock), .in1(_99));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4978 (.out1(R4979), .clock(clock), .in1(_59));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4979 (.out1(R4980), .clock(clock), .in1(_40));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op24 (.out1(_20), .in1(R4211));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op64 (.out1(_60), .in1(R4979), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op45 (.out1(_41), .in1(R4980), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op104 (.out1(_100), .in1(R4978), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op65 (.out1(_61), .in1(_41), .in2(_60));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op25 (.out1(_21), .in1(_20), .in2(2 'd 2));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op105 (.out1(_101), .in1(_61), .in2(_100));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op106 (.out1(_102), .in1(_101), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3700 (.out1(R3701), .clock(clock), .in1(R3700));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3956 (.out1(R3957), .clock(clock), .in1(R3956));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4211 (.out1(R4212), .clock(clock), .in1(R4211));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4456 (.out1(R4457), .clock(clock), .in1(R4456));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4696 (.out1(R4697), .clock(clock), .in1(R4696));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4980 (.out1(R4981), .clock(clock), .in1(_21));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4981 (.out1(R4982), .clock(clock), .in1(_102));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op107 (.out1(_103), .in1(R4982), .in2(57 'd 72340172838076673));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op26 (.out1(_22), .in1(base0_16_3544_D), .in2(R4981));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3701 (.out1(R3702), .clock(clock), .in1(R3701));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3957 (.out1(R3958), .clock(clock), .in1(R3957));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4212 (.out1(R4213), .clock(clock), .in1(R4212));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4457 (.out1(R4458), .clock(clock), .in1(R4457));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4697 (.out1(R4698), .clock(clock), .in1(R4697));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4982 (.out1(R4983), .clock(clock), .in1(_103));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4983 (.out1(R4984), .clock(clock), .in1(_22));
  SRAM op27 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_23),.ADR(R4984));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op108 (.out1(_104), .in1(R4983), .in2(6 'd 56));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3702 (.out1(R3703), .clock(clock), .in1(R3702));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3958 (.out1(R3959), .clock(clock), .in1(R3958));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4213 (.out1(R4214), .clock(clock), .in1(R4213));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4458 (.out1(R4459), .clock(clock), .in1(R4458));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4698 (.out1(R4699), .clock(clock), .in1(R4698));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4984 (.out1(R4985), .clock(clock), .in1(_23));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op4985 (.out1(R4986), .clock(clock), .in1(_104));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op109 (.out1(_105), .in1(R4986));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op110 (.out1(_106), .in1(R4985), .in2(_105));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op111 (.out1(idx_3545), .in1(_106), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3703 (.out1(R3704), .clock(clock), .in1(R3703));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3959 (.out1(R3960), .clock(clock), .in1(R3959));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4214 (.out1(R4215), .clock(clock), .in1(R4214));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4459 (.out1(R4460), .clock(clock), .in1(R4459));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4699 (.out1(R4700), .clock(clock), .in1(R4699));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4986 (.out1(R4987), .clock(clock), .in1(idx_3545));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op115 (.out1(_109), .in1(R4987));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op116 (.out1(_110), .in1(_109), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3704 (.out1(R3705), .clock(clock), .in1(R3704));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3960 (.out1(R3961), .clock(clock), .in1(R3960));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4215 (.out1(R4216), .clock(clock), .in1(R4215));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4460 (.out1(R4461), .clock(clock), .in1(R4460));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4700 (.out1(R4701), .clock(clock), .in1(R4700));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4987 (.out1(R4988), .clock(clock), .in1(R4987));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5219 (.out1(R5220), .clock(clock), .in1(_110));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op117 (.out1(_111), .in1(vec22_3547_D), .in2(R5220));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3705 (.out1(R3706), .clock(clock), .in1(R3705));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3961 (.out1(R3962), .clock(clock), .in1(R3961));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4216 (.out1(R4217), .clock(clock), .in1(R4216));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4461 (.out1(R4462), .clock(clock), .in1(R4461));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4701 (.out1(R4702), .clock(clock), .in1(R4701));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4988 (.out1(R4989), .clock(clock), .in1(R4988));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5220 (.out1(R5221), .clock(clock), .in1(_111));
  SRAM op118 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_112),.ADR(R5221));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3706 (.out1(R3707), .clock(clock), .in1(R3706));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3962 (.out1(R3963), .clock(clock), .in1(R3962));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4217 (.out1(R4218), .clock(clock), .in1(R4217));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4462 (.out1(R4463), .clock(clock), .in1(R4462));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4702 (.out1(R4703), .clock(clock), .in1(R4702));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4989 (.out1(R4990), .clock(clock), .in1(R4989));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5221 (.out1(R5222), .clock(clock), .in1(_112));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op112 (.out1(_107), .in1(ip1_3530_D), .in2(6 'd 36));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op113 (.out1(_108), .in1(_107));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op114 (.out1(off_3546), .in1(_108), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op119 (.out1(_113), .in1(R5222), .in2(off_3546));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3707 (.out1(R3708), .clock(clock), .in1(R3707));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3963 (.out1(R3964), .clock(clock), .in1(R3963));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4218 (.out1(R4219), .clock(clock), .in1(R4218));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4463 (.out1(R4464), .clock(clock), .in1(R4463));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4703 (.out1(R4704), .clock(clock), .in1(R4703));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4990 (.out1(R4991), .clock(clock), .in1(R4990));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5222 (.out1(R5223), .clock(clock), .in1(off_3546));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5449 (.out1(R5450), .clock(clock), .in1(_113));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op120 (.out1(_114), .in1(R5450), .in2(1 'd 1));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op121 (.out1(ifout121), .in1(_114), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op189 (.out1(_182), .in1(R4991));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op182 (.out1(_175), .in1(R4991));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op171 (.out1(_164), .in1(R4991));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op151 (.out1(_144), .in1(R4991));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op190 (.out1(_183), .in1(_182), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op183 (.out1(_176), .in1(_175), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op172 (.out1(_165), .in1(_164), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op152 (.out1(_145), .in1(_144), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3708 (.out1(R3709), .clock(clock), .in1(R3708));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3964 (.out1(R3965), .clock(clock), .in1(R3964));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4219 (.out1(R4220), .clock(clock), .in1(R4219));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4464 (.out1(R4465), .clock(clock), .in1(R4464));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4704 (.out1(R4705), .clock(clock), .in1(R4704));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4991 (.out1(R4992), .clock(clock), .in1(R4991));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5223 (.out1(R5224), .clock(clock), .in1(R5223));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5450 (.out1(R5451), .clock(clock), .in1(ifout121));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5684 (.out1(R5685), .clock(clock), .in1(_183));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5685 (.out1(R5686), .clock(clock), .in1(_176));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5686 (.out1(R5687), .clock(clock), .in1(_165));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5687 (.out1(R5688), .clock(clock), .in1(_145));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op164 (.out1(_157), .in1(R4992));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op144 (.out1(_137), .in1(R4992));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op133 (.out1(_126), .in1(R4992));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op126 (.out1(_119), .in1(R4992));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op193 (.out1(_186), .in1(2 'd 2), .in2(R5224));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op165 (.out1(_158), .in1(_157), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op145 (.out1(_138), .in1(_137), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op134 (.out1(_127), .in1(_126), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op127 (.out1(_120), .in1(_119), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op191 (.out1(_184), .in1(vec22_3547_D), .in2(R5685));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op184 (.out1(_177), .in1(vec22_3547_D), .in2(R5686));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op173 (.out1(_166), .in1(vec22_3547_D), .in2(R5687));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op153 (.out1(_146), .in1(vec22_3547_D), .in2(R5688));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3709 (.out1(R3710), .clock(clock), .in1(R3709));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3965 (.out1(R3966), .clock(clock), .in1(R3965));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4220 (.out1(R4221), .clock(clock), .in1(R4220));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4465 (.out1(R4466), .clock(clock), .in1(R4465));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4705 (.out1(R4706), .clock(clock), .in1(R4705));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4992 (.out1(R4993), .clock(clock), .in1(R4992));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5224 (.out1(R5225), .clock(clock), .in1(R5224));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5451 (.out1(R5452), .clock(clock), .in1(R5451));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5688 (.out1(R5689), .clock(clock), .in1(_186));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5689 (.out1(R5690), .clock(clock), .in1(_158));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5690 (.out1(R5691), .clock(clock), .in1(_138));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5691 (.out1(R5692), .clock(clock), .in1(_127));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5692 (.out1(R5693), .clock(clock), .in1(_120));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5693 (.out1(R5694), .clock(clock), .in1(_184));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5694 (.out1(R5695), .clock(clock), .in1(_177));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5695 (.out1(R5696), .clock(clock), .in1(_166));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5696 (.out1(R5697), .clock(clock), .in1(_146));
  SRAM op192 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_185),.ADR(R5694));
  SRAM op185 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_178),.ADR(R5695));
  SRAM op174 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_167),.ADR(R5696));
  SRAM op154 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_147),.ADR(R5697));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op186 (.out1(_179), .in1(2 'd 2), .in2(R5225));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op175 (.out1(_168), .in1(2 'd 2), .in2(R5225));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op168 (.out1(_161), .in1(2 'd 2), .in2(R5225));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op155 (.out1(_148), .in1(2 'd 2), .in2(R5225));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op148 (.out1(_141), .in1(2 'd 2), .in2(R5225));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op137 (.out1(_130), .in1(2 'd 2), .in2(R5225));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op166 (.out1(_159), .in1(vec22_3547_D), .in2(R5690));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op146 (.out1(_139), .in1(vec22_3547_D), .in2(R5691));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op135 (.out1(_128), .in1(vec22_3547_D), .in2(R5692));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op128 (.out1(_121), .in1(vec22_3547_D), .in2(R5693));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op194 (.out1(_187), .in1(R5689), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3710 (.out1(R3711), .clock(clock), .in1(R3710));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3966 (.out1(R3967), .clock(clock), .in1(R3966));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4221 (.out1(R4222), .clock(clock), .in1(R4221));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4466 (.out1(R4467), .clock(clock), .in1(R4466));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4706 (.out1(R4707), .clock(clock), .in1(R4706));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4993 (.out1(R4994), .clock(clock), .in1(R4993));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5225 (.out1(R5226), .clock(clock), .in1(R5225));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5452 (.out1(R5453), .clock(clock), .in1(R5452));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5697 (.out1(R5698), .clock(clock), .in1(_185));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5698 (.out1(R5699), .clock(clock), .in1(_178));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5699 (.out1(R5700), .clock(clock), .in1(_167));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5700 (.out1(R5701), .clock(clock), .in1(_147));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5701 (.out1(R5702), .clock(clock), .in1(_179));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5702 (.out1(R5703), .clock(clock), .in1(_168));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5703 (.out1(R5704), .clock(clock), .in1(_161));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5704 (.out1(R5705), .clock(clock), .in1(_148));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5705 (.out1(R5706), .clock(clock), .in1(_141));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5706 (.out1(R5707), .clock(clock), .in1(_130));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5707 (.out1(R5708), .clock(clock), .in1(_159));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5708 (.out1(R5709), .clock(clock), .in1(_139));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5709 (.out1(R5710), .clock(clock), .in1(_128));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5710 (.out1(R5711), .clock(clock), .in1(_121));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5711 (.out1(R5712), .clock(clock), .in1(_187));
  SRAM op167 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_160),.ADR(R5708));
  SRAM op147 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_140),.ADR(R5709));
  SRAM op136 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_129),.ADR(R5710));
  SRAM op129 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_122),.ADR(R5711));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op195 (.out1(_188), .in1(R5698), .in2(R5712));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op196 (.out1(_189), .in1(_188), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op187 (.out1(_180), .in1(R5702), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op176 (.out1(_169), .in1(R5703), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op156 (.out1(_149), .in1(R5705), .in2(64 'd 18446744073709551615));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op130 (.out1(_123), .in1(2 'd 2), .in2(R5226));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op197 (.out1(_190), .in1(_189), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op188 (.out1(_181), .in1(R5699), .in2(_180));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op177 (.out1(_170), .in1(R5700), .in2(_169));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op157 (.out1(_150), .in1(R5701), .in2(_149));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op198 (.out1(_191), .in1(_181), .in2(_190));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op178 (.out1(_171), .in1(_170), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op169 (.out1(_162), .in1(R5704), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op158 (.out1(_151), .in1(_150), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op149 (.out1(_142), .in1(R5706), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op138 (.out1(_131), .in1(R5707), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3711 (.out1(R3712), .clock(clock), .in1(R3711));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3967 (.out1(R3968), .clock(clock), .in1(R3967));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4222 (.out1(R4223), .clock(clock), .in1(R4222));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4467 (.out1(R4468), .clock(clock), .in1(R4467));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4707 (.out1(R4708), .clock(clock), .in1(R4707));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4994 (.out1(R4995), .clock(clock), .in1(R4994));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5226 (.out1(R5227), .clock(clock), .in1(R5226));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5453 (.out1(R5454), .clock(clock), .in1(R5453));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5712 (.out1(R5713), .clock(clock), .in1(_160));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5713 (.out1(R5714), .clock(clock), .in1(_140));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5714 (.out1(R5715), .clock(clock), .in1(_129));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5715 (.out1(R5716), .clock(clock), .in1(_122));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5716 (.out1(R5717), .clock(clock), .in1(_123));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5717 (.out1(R5718), .clock(clock), .in1(_191));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5718 (.out1(R5719), .clock(clock), .in1(_171));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5719 (.out1(R5720), .clock(clock), .in1(_162));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5720 (.out1(R5721), .clock(clock), .in1(_151));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5721 (.out1(R5722), .clock(clock), .in1(_142));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5722 (.out1(R5723), .clock(clock), .in1(_131));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op179 (.out1(_172), .in1(R5719), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op170 (.out1(_163), .in1(R5713), .in2(R5720));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op139 (.out1(_132), .in1(R5715), .in2(R5723));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op199 (.out1(_192), .in1(R5718), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op180 (.out1(_173), .in1(_163), .in2(_172));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op159 (.out1(_152), .in1(R5721), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op150 (.out1(_143), .in1(R5714), .in2(R5722));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op140 (.out1(_133), .in1(_132), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op131 (.out1(_124), .in1(R5717), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op160 (.out1(_153), .in1(_143), .in2(_152));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op200 (.out1(_193), .in1(_192), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op181 (.out1(_174), .in1(_173), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op141 (.out1(_134), .in1(_133), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op132 (.out1(_125), .in1(R5716), .in2(_124));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op201 (.out1(_194), .in1(_174), .in2(_193));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op161 (.out1(_154), .in1(_153), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op142 (.out1(_135), .in1(_125), .in2(_134));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3712 (.out1(R3713), .clock(clock), .in1(R3712));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3968 (.out1(R3969), .clock(clock), .in1(R3968));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4223 (.out1(R4224), .clock(clock), .in1(R4223));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4468 (.out1(R4469), .clock(clock), .in1(R4468));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4708 (.out1(R4709), .clock(clock), .in1(R4708));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4995 (.out1(R4996), .clock(clock), .in1(R4995));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5227 (.out1(R5228), .clock(clock), .in1(R5227));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5454 (.out1(R5455), .clock(clock), .in1(R5454));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5723 (.out1(R5724), .clock(clock), .in1(_194));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5724 (.out1(R5725), .clock(clock), .in1(_154));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5725 (.out1(R5726), .clock(clock), .in1(_135));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op122 (.out1(_115), .in1(R4996));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op162 (.out1(_155), .in1(R5725), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op143 (.out1(_136), .in1(R5726), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op202 (.out1(_195), .in1(R5724), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op163 (.out1(_156), .in1(_136), .in2(_155));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op123 (.out1(_116), .in1(_115), .in2(2 'd 2));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op203 (.out1(_196), .in1(_156), .in2(_195));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op204 (.out1(_197), .in1(_196), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3713 (.out1(R3714), .clock(clock), .in1(R3713));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3969 (.out1(R3970), .clock(clock), .in1(R3969));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4224 (.out1(R4225), .clock(clock), .in1(R4224));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4469 (.out1(R4470), .clock(clock), .in1(R4469));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4709 (.out1(R4710), .clock(clock), .in1(R4709));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4996 (.out1(R4997), .clock(clock), .in1(R4996));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5228 (.out1(R5229), .clock(clock), .in1(R5228));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5455 (.out1(R5456), .clock(clock), .in1(R5455));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5726 (.out1(R5727), .clock(clock), .in1(_116));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5727 (.out1(R5728), .clock(clock), .in1(_197));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op205 (.out1(_198), .in1(R5728), .in2(57 'd 72340172838076673));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op124 (.out1(_117), .in1(base0_22_3552_D), .in2(R5727));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3714 (.out1(R3715), .clock(clock), .in1(R3714));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3970 (.out1(R3971), .clock(clock), .in1(R3970));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4225 (.out1(R4226), .clock(clock), .in1(R4225));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4470 (.out1(R4471), .clock(clock), .in1(R4470));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4710 (.out1(R4711), .clock(clock), .in1(R4710));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4997 (.out1(R4998), .clock(clock), .in1(R4997));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5229 (.out1(R5230), .clock(clock), .in1(R5229));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5456 (.out1(R5457), .clock(clock), .in1(R5456));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5728 (.out1(R5729), .clock(clock), .in1(_198));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5729 (.out1(R5730), .clock(clock), .in1(_117));
  SRAM op125 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_118),.ADR(R5730));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op206 (.out1(_199), .in1(R5729), .in2(6 'd 56));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3715 (.out1(R3716), .clock(clock), .in1(R3715));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3971 (.out1(R3972), .clock(clock), .in1(R3971));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4226 (.out1(R4227), .clock(clock), .in1(R4226));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4471 (.out1(R4472), .clock(clock), .in1(R4471));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4711 (.out1(R4712), .clock(clock), .in1(R4711));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4998 (.out1(R4999), .clock(clock), .in1(R4998));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5230 (.out1(R5231), .clock(clock), .in1(R5230));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5457 (.out1(R5458), .clock(clock), .in1(R5457));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5730 (.out1(R5731), .clock(clock), .in1(_118));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5731 (.out1(R5732), .clock(clock), .in1(_199));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op207 (.out1(_200), .in1(R5732));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op208 (.out1(_201), .in1(R5731), .in2(_200));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op209 (.out1(idx_3553), .in1(_201), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3716 (.out1(R3717), .clock(clock), .in1(R3716));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3972 (.out1(R3973), .clock(clock), .in1(R3972));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4227 (.out1(R4228), .clock(clock), .in1(R4227));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4472 (.out1(R4473), .clock(clock), .in1(R4472));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4712 (.out1(R4713), .clock(clock), .in1(R4712));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4999 (.out1(R5000), .clock(clock), .in1(R4999));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5231 (.out1(R5232), .clock(clock), .in1(R5231));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5458 (.out1(R5459), .clock(clock), .in1(R5458));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5732 (.out1(R5733), .clock(clock), .in1(idx_3553));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op213 (.out1(_204), .in1(R5733));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op214 (.out1(_205), .in1(_204), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3717 (.out1(R3718), .clock(clock), .in1(R3717));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3973 (.out1(R3974), .clock(clock), .in1(R3973));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4228 (.out1(R4229), .clock(clock), .in1(R4228));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4473 (.out1(R4474), .clock(clock), .in1(R4473));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4713 (.out1(R4714), .clock(clock), .in1(R4713));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5000 (.out1(R5001), .clock(clock), .in1(R5000));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5232 (.out1(R5233), .clock(clock), .in1(R5232));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5459 (.out1(R5460), .clock(clock), .in1(R5459));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5733 (.out1(R5734), .clock(clock), .in1(R5733));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5951 (.out1(R5952), .clock(clock), .in1(_205));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op215 (.out1(_206), .in1(vec28_3555_D), .in2(R5952));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3718 (.out1(R3719), .clock(clock), .in1(R3718));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3974 (.out1(R3975), .clock(clock), .in1(R3974));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4229 (.out1(R4230), .clock(clock), .in1(R4229));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4474 (.out1(R4475), .clock(clock), .in1(R4474));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4714 (.out1(R4715), .clock(clock), .in1(R4714));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5001 (.out1(R5002), .clock(clock), .in1(R5001));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5233 (.out1(R5234), .clock(clock), .in1(R5233));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5460 (.out1(R5461), .clock(clock), .in1(R5460));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5734 (.out1(R5735), .clock(clock), .in1(R5734));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5952 (.out1(R5953), .clock(clock), .in1(_206));
  SRAM op216 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_207),.ADR(R5953));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3719 (.out1(R3720), .clock(clock), .in1(R3719));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3975 (.out1(R3976), .clock(clock), .in1(R3975));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4230 (.out1(R4231), .clock(clock), .in1(R4230));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4475 (.out1(R4476), .clock(clock), .in1(R4475));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4715 (.out1(R4716), .clock(clock), .in1(R4715));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5002 (.out1(R5003), .clock(clock), .in1(R5002));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5234 (.out1(R5235), .clock(clock), .in1(R5234));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5461 (.out1(R5462), .clock(clock), .in1(R5461));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5735 (.out1(R5736), .clock(clock), .in1(R5735));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op5953 (.out1(R5954), .clock(clock), .in1(_207));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(5), .BITSIZE_out1(64), .PRECISION(64)) op210 (.out1(_202), .in1(ip1_3530_D), .in2(5 'd 30));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op211 (.out1(_203), .in1(_202));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op212 (.out1(off_3554), .in1(_203), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op217 (.out1(_208), .in1(R5954), .in2(off_3554));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3720 (.out1(R3721), .clock(clock), .in1(R3720));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3976 (.out1(R3977), .clock(clock), .in1(R3976));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4231 (.out1(R4232), .clock(clock), .in1(R4231));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4476 (.out1(R4477), .clock(clock), .in1(R4476));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4716 (.out1(R4717), .clock(clock), .in1(R4716));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5003 (.out1(R5004), .clock(clock), .in1(R5003));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5235 (.out1(R5236), .clock(clock), .in1(R5235));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5462 (.out1(R5463), .clock(clock), .in1(R5462));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5736 (.out1(R5737), .clock(clock), .in1(R5736));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5954 (.out1(R5955), .clock(clock), .in1(off_3554));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6167 (.out1(R6168), .clock(clock), .in1(_208));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op218 (.out1(_209), .in1(R6168), .in2(1 'd 1));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op219 (.out1(ifout219), .in1(_209), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op287 (.out1(_277), .in1(R5737));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op280 (.out1(_270), .in1(R5737));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op269 (.out1(_259), .in1(R5737));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op249 (.out1(_239), .in1(R5737));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op288 (.out1(_278), .in1(_277), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op281 (.out1(_271), .in1(_270), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op270 (.out1(_260), .in1(_259), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op250 (.out1(_240), .in1(_239), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3721 (.out1(R3722), .clock(clock), .in1(R3721));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3977 (.out1(R3978), .clock(clock), .in1(R3977));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4232 (.out1(R4233), .clock(clock), .in1(R4232));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4477 (.out1(R4478), .clock(clock), .in1(R4477));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4717 (.out1(R4718), .clock(clock), .in1(R4717));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5004 (.out1(R5005), .clock(clock), .in1(R5004));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5236 (.out1(R5237), .clock(clock), .in1(R5236));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5463 (.out1(R5464), .clock(clock), .in1(R5463));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5737 (.out1(R5738), .clock(clock), .in1(R5737));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5955 (.out1(R5956), .clock(clock), .in1(R5955));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6168 (.out1(R6169), .clock(clock), .in1(ifout219));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6389 (.out1(R6390), .clock(clock), .in1(_278));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6390 (.out1(R6391), .clock(clock), .in1(_271));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6391 (.out1(R6392), .clock(clock), .in1(_260));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6392 (.out1(R6393), .clock(clock), .in1(_240));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op262 (.out1(_252), .in1(R5738));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op242 (.out1(_232), .in1(R5738));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op231 (.out1(_221), .in1(R5738));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op224 (.out1(_214), .in1(R5738));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op291 (.out1(_281), .in1(2 'd 2), .in2(R5956));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op263 (.out1(_253), .in1(_252), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op243 (.out1(_233), .in1(_232), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op232 (.out1(_222), .in1(_221), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op225 (.out1(_215), .in1(_214), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op289 (.out1(_279), .in1(vec28_3555_D), .in2(R6390));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op282 (.out1(_272), .in1(vec28_3555_D), .in2(R6391));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op271 (.out1(_261), .in1(vec28_3555_D), .in2(R6392));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op251 (.out1(_241), .in1(vec28_3555_D), .in2(R6393));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3722 (.out1(R3723), .clock(clock), .in1(R3722));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3978 (.out1(R3979), .clock(clock), .in1(R3978));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4233 (.out1(R4234), .clock(clock), .in1(R4233));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4478 (.out1(R4479), .clock(clock), .in1(R4478));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4718 (.out1(R4719), .clock(clock), .in1(R4718));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5005 (.out1(R5006), .clock(clock), .in1(R5005));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5237 (.out1(R5238), .clock(clock), .in1(R5237));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5464 (.out1(R5465), .clock(clock), .in1(R5464));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5738 (.out1(R5739), .clock(clock), .in1(R5738));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5956 (.out1(R5957), .clock(clock), .in1(R5956));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6169 (.out1(R6170), .clock(clock), .in1(R6169));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6393 (.out1(R6394), .clock(clock), .in1(_281));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6394 (.out1(R6395), .clock(clock), .in1(_253));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6395 (.out1(R6396), .clock(clock), .in1(_233));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6396 (.out1(R6397), .clock(clock), .in1(_222));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6397 (.out1(R6398), .clock(clock), .in1(_215));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6398 (.out1(R6399), .clock(clock), .in1(_279));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6399 (.out1(R6400), .clock(clock), .in1(_272));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6400 (.out1(R6401), .clock(clock), .in1(_261));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6401 (.out1(R6402), .clock(clock), .in1(_241));
  SRAM op290 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_280),.ADR(R6399));
  SRAM op283 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_273),.ADR(R6400));
  SRAM op272 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_262),.ADR(R6401));
  SRAM op252 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_242),.ADR(R6402));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op284 (.out1(_274), .in1(2 'd 2), .in2(R5957));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op273 (.out1(_263), .in1(2 'd 2), .in2(R5957));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op266 (.out1(_256), .in1(2 'd 2), .in2(R5957));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op253 (.out1(_243), .in1(2 'd 2), .in2(R5957));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op246 (.out1(_236), .in1(2 'd 2), .in2(R5957));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op235 (.out1(_225), .in1(2 'd 2), .in2(R5957));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op264 (.out1(_254), .in1(vec28_3555_D), .in2(R6395));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op244 (.out1(_234), .in1(vec28_3555_D), .in2(R6396));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op233 (.out1(_223), .in1(vec28_3555_D), .in2(R6397));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op226 (.out1(_216), .in1(vec28_3555_D), .in2(R6398));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op292 (.out1(_282), .in1(R6394), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3723 (.out1(R3724), .clock(clock), .in1(R3723));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3979 (.out1(R3980), .clock(clock), .in1(R3979));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4234 (.out1(R4235), .clock(clock), .in1(R4234));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4479 (.out1(R4480), .clock(clock), .in1(R4479));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4719 (.out1(R4720), .clock(clock), .in1(R4719));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5006 (.out1(R5007), .clock(clock), .in1(R5006));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5238 (.out1(R5239), .clock(clock), .in1(R5238));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5465 (.out1(R5466), .clock(clock), .in1(R5465));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5739 (.out1(R5740), .clock(clock), .in1(R5739));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5957 (.out1(R5958), .clock(clock), .in1(R5957));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6170 (.out1(R6171), .clock(clock), .in1(R6170));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6402 (.out1(R6403), .clock(clock), .in1(_280));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6403 (.out1(R6404), .clock(clock), .in1(_273));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6404 (.out1(R6405), .clock(clock), .in1(_262));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6405 (.out1(R6406), .clock(clock), .in1(_242));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6406 (.out1(R6407), .clock(clock), .in1(_274));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6407 (.out1(R6408), .clock(clock), .in1(_263));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6408 (.out1(R6409), .clock(clock), .in1(_256));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6409 (.out1(R6410), .clock(clock), .in1(_243));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6410 (.out1(R6411), .clock(clock), .in1(_236));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6411 (.out1(R6412), .clock(clock), .in1(_225));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6412 (.out1(R6413), .clock(clock), .in1(_254));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6413 (.out1(R6414), .clock(clock), .in1(_234));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6414 (.out1(R6415), .clock(clock), .in1(_223));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6415 (.out1(R6416), .clock(clock), .in1(_216));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6416 (.out1(R6417), .clock(clock), .in1(_282));
  SRAM op265 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_255),.ADR(R6413));
  SRAM op245 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_235),.ADR(R6414));
  SRAM op234 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_224),.ADR(R6415));
  SRAM op227 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_217),.ADR(R6416));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op293 (.out1(_283), .in1(R6403), .in2(R6417));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op294 (.out1(_284), .in1(_283), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op285 (.out1(_275), .in1(R6407), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op274 (.out1(_264), .in1(R6408), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op254 (.out1(_244), .in1(R6410), .in2(64 'd 18446744073709551615));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op228 (.out1(_218), .in1(2 'd 2), .in2(R5958));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op295 (.out1(_285), .in1(_284), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op286 (.out1(_276), .in1(R6404), .in2(_275));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op275 (.out1(_265), .in1(R6405), .in2(_264));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op255 (.out1(_245), .in1(R6406), .in2(_244));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op296 (.out1(_286), .in1(_276), .in2(_285));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op276 (.out1(_266), .in1(_265), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op267 (.out1(_257), .in1(R6409), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op256 (.out1(_246), .in1(_245), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op247 (.out1(_237), .in1(R6411), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op236 (.out1(_226), .in1(R6412), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3724 (.out1(R3725), .clock(clock), .in1(R3724));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3980 (.out1(R3981), .clock(clock), .in1(R3980));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4235 (.out1(R4236), .clock(clock), .in1(R4235));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4480 (.out1(R4481), .clock(clock), .in1(R4480));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4720 (.out1(R4721), .clock(clock), .in1(R4720));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5007 (.out1(R5008), .clock(clock), .in1(R5007));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5239 (.out1(R5240), .clock(clock), .in1(R5239));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5466 (.out1(R5467), .clock(clock), .in1(R5466));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5740 (.out1(R5741), .clock(clock), .in1(R5740));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5958 (.out1(R5959), .clock(clock), .in1(R5958));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6171 (.out1(R6172), .clock(clock), .in1(R6171));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6417 (.out1(R6418), .clock(clock), .in1(_255));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6418 (.out1(R6419), .clock(clock), .in1(_235));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6419 (.out1(R6420), .clock(clock), .in1(_224));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6420 (.out1(R6421), .clock(clock), .in1(_217));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6421 (.out1(R6422), .clock(clock), .in1(_218));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6422 (.out1(R6423), .clock(clock), .in1(_286));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6423 (.out1(R6424), .clock(clock), .in1(_266));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6424 (.out1(R6425), .clock(clock), .in1(_257));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6425 (.out1(R6426), .clock(clock), .in1(_246));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6426 (.out1(R6427), .clock(clock), .in1(_237));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6427 (.out1(R6428), .clock(clock), .in1(_226));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op277 (.out1(_267), .in1(R6424), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op268 (.out1(_258), .in1(R6418), .in2(R6425));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op237 (.out1(_227), .in1(R6420), .in2(R6428));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op297 (.out1(_287), .in1(R6423), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op278 (.out1(_268), .in1(_258), .in2(_267));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op257 (.out1(_247), .in1(R6426), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op248 (.out1(_238), .in1(R6419), .in2(R6427));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op238 (.out1(_228), .in1(_227), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op229 (.out1(_219), .in1(R6422), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op258 (.out1(_248), .in1(_238), .in2(_247));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op298 (.out1(_288), .in1(_287), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op279 (.out1(_269), .in1(_268), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op239 (.out1(_229), .in1(_228), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op230 (.out1(_220), .in1(R6421), .in2(_219));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op299 (.out1(_289), .in1(_269), .in2(_288));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op259 (.out1(_249), .in1(_248), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op240 (.out1(_230), .in1(_220), .in2(_229));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3725 (.out1(R3726), .clock(clock), .in1(R3725));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3981 (.out1(R3982), .clock(clock), .in1(R3981));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4236 (.out1(R4237), .clock(clock), .in1(R4236));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4481 (.out1(R4482), .clock(clock), .in1(R4481));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4721 (.out1(R4722), .clock(clock), .in1(R4721));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5008 (.out1(R5009), .clock(clock), .in1(R5008));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5240 (.out1(R5241), .clock(clock), .in1(R5240));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5467 (.out1(R5468), .clock(clock), .in1(R5467));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5741 (.out1(R5742), .clock(clock), .in1(R5741));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5959 (.out1(R5960), .clock(clock), .in1(R5959));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6172 (.out1(R6173), .clock(clock), .in1(R6172));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6428 (.out1(R6429), .clock(clock), .in1(_289));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6429 (.out1(R6430), .clock(clock), .in1(_249));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6430 (.out1(R6431), .clock(clock), .in1(_230));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op220 (.out1(_210), .in1(R5742));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op260 (.out1(_250), .in1(R6430), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op241 (.out1(_231), .in1(R6431), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op300 (.out1(_290), .in1(R6429), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op261 (.out1(_251), .in1(_231), .in2(_250));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op221 (.out1(_211), .in1(_210), .in2(2 'd 2));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op301 (.out1(_291), .in1(_251), .in2(_290));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op302 (.out1(_292), .in1(_291), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3726 (.out1(R3727), .clock(clock), .in1(R3726));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3982 (.out1(R3983), .clock(clock), .in1(R3982));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4237 (.out1(R4238), .clock(clock), .in1(R4237));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4482 (.out1(R4483), .clock(clock), .in1(R4482));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4722 (.out1(R4723), .clock(clock), .in1(R4722));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5009 (.out1(R5010), .clock(clock), .in1(R5009));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5241 (.out1(R5242), .clock(clock), .in1(R5241));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5468 (.out1(R5469), .clock(clock), .in1(R5468));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5742 (.out1(R5743), .clock(clock), .in1(R5742));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5960 (.out1(R5961), .clock(clock), .in1(R5960));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6173 (.out1(R6174), .clock(clock), .in1(R6173));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6431 (.out1(R6432), .clock(clock), .in1(_211));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6432 (.out1(R6433), .clock(clock), .in1(_292));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op303 (.out1(_293), .in1(R6433), .in2(57 'd 72340172838076673));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op222 (.out1(_212), .in1(base0_28_3560_D), .in2(R6432));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3727 (.out1(R3728), .clock(clock), .in1(R3727));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3983 (.out1(R3984), .clock(clock), .in1(R3983));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4238 (.out1(R4239), .clock(clock), .in1(R4238));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4483 (.out1(R4484), .clock(clock), .in1(R4483));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4723 (.out1(R4724), .clock(clock), .in1(R4723));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5010 (.out1(R5011), .clock(clock), .in1(R5010));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5242 (.out1(R5243), .clock(clock), .in1(R5242));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5469 (.out1(R5470), .clock(clock), .in1(R5469));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5743 (.out1(R5744), .clock(clock), .in1(R5743));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5961 (.out1(R5962), .clock(clock), .in1(R5961));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6174 (.out1(R6175), .clock(clock), .in1(R6174));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6433 (.out1(R6434), .clock(clock), .in1(_293));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6434 (.out1(R6435), .clock(clock), .in1(_212));
  SRAM op223 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_213),.ADR(R6435));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op304 (.out1(_294), .in1(R6434), .in2(6 'd 56));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3728 (.out1(R3729), .clock(clock), .in1(R3728));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3984 (.out1(R3985), .clock(clock), .in1(R3984));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4239 (.out1(R4240), .clock(clock), .in1(R4239));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4484 (.out1(R4485), .clock(clock), .in1(R4484));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4724 (.out1(R4725), .clock(clock), .in1(R4724));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5011 (.out1(R5012), .clock(clock), .in1(R5011));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5243 (.out1(R5244), .clock(clock), .in1(R5243));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5470 (.out1(R5471), .clock(clock), .in1(R5470));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5744 (.out1(R5745), .clock(clock), .in1(R5744));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5962 (.out1(R5963), .clock(clock), .in1(R5962));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6175 (.out1(R6176), .clock(clock), .in1(R6175));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6435 (.out1(R6436), .clock(clock), .in1(_213));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6436 (.out1(R6437), .clock(clock), .in1(_294));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op305 (.out1(_295), .in1(R6437));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op306 (.out1(_296), .in1(R6436), .in2(_295));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op307 (.out1(idx_3561), .in1(_296), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3729 (.out1(R3730), .clock(clock), .in1(R3729));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3985 (.out1(R3986), .clock(clock), .in1(R3985));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4240 (.out1(R4241), .clock(clock), .in1(R4240));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4485 (.out1(R4486), .clock(clock), .in1(R4485));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4725 (.out1(R4726), .clock(clock), .in1(R4725));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5012 (.out1(R5013), .clock(clock), .in1(R5012));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5244 (.out1(R5245), .clock(clock), .in1(R5244));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5471 (.out1(R5472), .clock(clock), .in1(R5471));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5745 (.out1(R5746), .clock(clock), .in1(R5745));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5963 (.out1(R5964), .clock(clock), .in1(R5963));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6176 (.out1(R6177), .clock(clock), .in1(R6176));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6437 (.out1(R6438), .clock(clock), .in1(idx_3561));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op311 (.out1(_299), .in1(R6438));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op312 (.out1(_300), .in1(_299), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3730 (.out1(R3731), .clock(clock), .in1(R3730));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3986 (.out1(R3987), .clock(clock), .in1(R3986));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4241 (.out1(R4242), .clock(clock), .in1(R4241));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4486 (.out1(R4487), .clock(clock), .in1(R4486));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4726 (.out1(R4727), .clock(clock), .in1(R4726));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5013 (.out1(R5014), .clock(clock), .in1(R5013));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5245 (.out1(R5246), .clock(clock), .in1(R5245));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5472 (.out1(R5473), .clock(clock), .in1(R5472));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5746 (.out1(R5747), .clock(clock), .in1(R5746));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5964 (.out1(R5965), .clock(clock), .in1(R5964));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6177 (.out1(R6178), .clock(clock), .in1(R6177));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6438 (.out1(R6439), .clock(clock), .in1(R6438));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6643 (.out1(R6644), .clock(clock), .in1(_300));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op313 (.out1(_301), .in1(vec34_3563_D), .in2(R6644));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3731 (.out1(R3732), .clock(clock), .in1(R3731));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3987 (.out1(R3988), .clock(clock), .in1(R3987));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4242 (.out1(R4243), .clock(clock), .in1(R4242));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4487 (.out1(R4488), .clock(clock), .in1(R4487));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4727 (.out1(R4728), .clock(clock), .in1(R4727));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5014 (.out1(R5015), .clock(clock), .in1(R5014));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5246 (.out1(R5247), .clock(clock), .in1(R5246));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5473 (.out1(R5474), .clock(clock), .in1(R5473));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5747 (.out1(R5748), .clock(clock), .in1(R5747));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5965 (.out1(R5966), .clock(clock), .in1(R5965));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6178 (.out1(R6179), .clock(clock), .in1(R6178));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6439 (.out1(R6440), .clock(clock), .in1(R6439));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6644 (.out1(R6645), .clock(clock), .in1(_301));
  SRAM op314 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_302),.ADR(R6645));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3732 (.out1(R3733), .clock(clock), .in1(R3732));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3988 (.out1(R3989), .clock(clock), .in1(R3988));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4243 (.out1(R4244), .clock(clock), .in1(R4243));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4488 (.out1(R4489), .clock(clock), .in1(R4488));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4728 (.out1(R4729), .clock(clock), .in1(R4728));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5015 (.out1(R5016), .clock(clock), .in1(R5015));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5247 (.out1(R5248), .clock(clock), .in1(R5247));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5474 (.out1(R5475), .clock(clock), .in1(R5474));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5748 (.out1(R5749), .clock(clock), .in1(R5748));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5966 (.out1(R5967), .clock(clock), .in1(R5966));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6179 (.out1(R6180), .clock(clock), .in1(R6179));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6440 (.out1(R6441), .clock(clock), .in1(R6440));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6645 (.out1(R6646), .clock(clock), .in1(_302));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(5), .BITSIZE_out1(64), .PRECISION(64)) op308 (.out1(_297), .in1(ip1_3530_D), .in2(5 'd 24));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op309 (.out1(_298), .in1(_297));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op310 (.out1(off_3562), .in1(_298), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op315 (.out1(_303), .in1(R6646), .in2(off_3562));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3733 (.out1(R3734), .clock(clock), .in1(R3733));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3989 (.out1(R3990), .clock(clock), .in1(R3989));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4244 (.out1(R4245), .clock(clock), .in1(R4244));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4489 (.out1(R4490), .clock(clock), .in1(R4489));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4729 (.out1(R4730), .clock(clock), .in1(R4729));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5016 (.out1(R5017), .clock(clock), .in1(R5016));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5248 (.out1(R5249), .clock(clock), .in1(R5248));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5475 (.out1(R5476), .clock(clock), .in1(R5475));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5749 (.out1(R5750), .clock(clock), .in1(R5749));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5967 (.out1(R5968), .clock(clock), .in1(R5967));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6180 (.out1(R6181), .clock(clock), .in1(R6180));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6441 (.out1(R6442), .clock(clock), .in1(R6441));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6646 (.out1(R6647), .clock(clock), .in1(off_3562));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op6846 (.out1(R6847), .clock(clock), .in1(_303));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op316 (.out1(_304), .in1(R6847), .in2(1 'd 1));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op317 (.out1(ifout317), .in1(_304), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op385 (.out1(_372), .in1(R6442));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op378 (.out1(_365), .in1(R6442));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op367 (.out1(_354), .in1(R6442));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op347 (.out1(_334), .in1(R6442));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op386 (.out1(_373), .in1(_372), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op379 (.out1(_366), .in1(_365), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op368 (.out1(_355), .in1(_354), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op348 (.out1(_335), .in1(_334), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3734 (.out1(R3735), .clock(clock), .in1(R3734));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3990 (.out1(R3991), .clock(clock), .in1(R3990));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4245 (.out1(R4246), .clock(clock), .in1(R4245));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4490 (.out1(R4491), .clock(clock), .in1(R4490));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4730 (.out1(R4731), .clock(clock), .in1(R4730));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5017 (.out1(R5018), .clock(clock), .in1(R5017));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5249 (.out1(R5250), .clock(clock), .in1(R5249));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5476 (.out1(R5477), .clock(clock), .in1(R5476));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5750 (.out1(R5751), .clock(clock), .in1(R5750));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5968 (.out1(R5969), .clock(clock), .in1(R5968));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6181 (.out1(R6182), .clock(clock), .in1(R6181));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6442 (.out1(R6443), .clock(clock), .in1(R6442));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6647 (.out1(R6648), .clock(clock), .in1(R6647));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6847 (.out1(R6848), .clock(clock), .in1(ifout317));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7054 (.out1(R7055), .clock(clock), .in1(_373));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7055 (.out1(R7056), .clock(clock), .in1(_366));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7056 (.out1(R7057), .clock(clock), .in1(_355));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7057 (.out1(R7058), .clock(clock), .in1(_335));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op360 (.out1(_347), .in1(R6443));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op340 (.out1(_327), .in1(R6443));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op329 (.out1(_316), .in1(R6443));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op322 (.out1(_309), .in1(R6443));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op389 (.out1(_376), .in1(2 'd 2), .in2(R6648));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op361 (.out1(_348), .in1(_347), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op341 (.out1(_328), .in1(_327), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op330 (.out1(_317), .in1(_316), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op323 (.out1(_310), .in1(_309), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op387 (.out1(_374), .in1(vec34_3563_D), .in2(R7055));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op380 (.out1(_367), .in1(vec34_3563_D), .in2(R7056));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op369 (.out1(_356), .in1(vec34_3563_D), .in2(R7057));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op349 (.out1(_336), .in1(vec34_3563_D), .in2(R7058));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3735 (.out1(R3736), .clock(clock), .in1(R3735));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3991 (.out1(R3992), .clock(clock), .in1(R3991));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4246 (.out1(R4247), .clock(clock), .in1(R4246));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4491 (.out1(R4492), .clock(clock), .in1(R4491));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4731 (.out1(R4732), .clock(clock), .in1(R4731));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5018 (.out1(R5019), .clock(clock), .in1(R5018));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5250 (.out1(R5251), .clock(clock), .in1(R5250));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5477 (.out1(R5478), .clock(clock), .in1(R5477));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5751 (.out1(R5752), .clock(clock), .in1(R5751));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5969 (.out1(R5970), .clock(clock), .in1(R5969));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6182 (.out1(R6183), .clock(clock), .in1(R6182));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6443 (.out1(R6444), .clock(clock), .in1(R6443));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6648 (.out1(R6649), .clock(clock), .in1(R6648));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6848 (.out1(R6849), .clock(clock), .in1(R6848));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7058 (.out1(R7059), .clock(clock), .in1(_376));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7059 (.out1(R7060), .clock(clock), .in1(_348));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7060 (.out1(R7061), .clock(clock), .in1(_328));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7061 (.out1(R7062), .clock(clock), .in1(_317));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7062 (.out1(R7063), .clock(clock), .in1(_310));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7063 (.out1(R7064), .clock(clock), .in1(_374));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7064 (.out1(R7065), .clock(clock), .in1(_367));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7065 (.out1(R7066), .clock(clock), .in1(_356));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7066 (.out1(R7067), .clock(clock), .in1(_336));
  SRAM op388 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_375),.ADR(R7064));
  SRAM op381 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_368),.ADR(R7065));
  SRAM op370 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_357),.ADR(R7066));
  SRAM op350 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_337),.ADR(R7067));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op382 (.out1(_369), .in1(2 'd 2), .in2(R6649));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op371 (.out1(_358), .in1(2 'd 2), .in2(R6649));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op364 (.out1(_351), .in1(2 'd 2), .in2(R6649));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op351 (.out1(_338), .in1(2 'd 2), .in2(R6649));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op344 (.out1(_331), .in1(2 'd 2), .in2(R6649));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op333 (.out1(_320), .in1(2 'd 2), .in2(R6649));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op362 (.out1(_349), .in1(vec34_3563_D), .in2(R7060));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op342 (.out1(_329), .in1(vec34_3563_D), .in2(R7061));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op331 (.out1(_318), .in1(vec34_3563_D), .in2(R7062));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op324 (.out1(_311), .in1(vec34_3563_D), .in2(R7063));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op390 (.out1(_377), .in1(R7059), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3736 (.out1(R3737), .clock(clock), .in1(R3736));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3992 (.out1(R3993), .clock(clock), .in1(R3992));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4247 (.out1(R4248), .clock(clock), .in1(R4247));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4492 (.out1(R4493), .clock(clock), .in1(R4492));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4732 (.out1(R4733), .clock(clock), .in1(R4732));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5019 (.out1(R5020), .clock(clock), .in1(R5019));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5251 (.out1(R5252), .clock(clock), .in1(R5251));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5478 (.out1(R5479), .clock(clock), .in1(R5478));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5752 (.out1(R5753), .clock(clock), .in1(R5752));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5970 (.out1(R5971), .clock(clock), .in1(R5970));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6183 (.out1(R6184), .clock(clock), .in1(R6183));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6444 (.out1(R6445), .clock(clock), .in1(R6444));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6649 (.out1(R6650), .clock(clock), .in1(R6649));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6849 (.out1(R6850), .clock(clock), .in1(R6849));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7067 (.out1(R7068), .clock(clock), .in1(_375));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7068 (.out1(R7069), .clock(clock), .in1(_368));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7069 (.out1(R7070), .clock(clock), .in1(_357));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7070 (.out1(R7071), .clock(clock), .in1(_337));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7071 (.out1(R7072), .clock(clock), .in1(_369));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7072 (.out1(R7073), .clock(clock), .in1(_358));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7073 (.out1(R7074), .clock(clock), .in1(_351));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7074 (.out1(R7075), .clock(clock), .in1(_338));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7075 (.out1(R7076), .clock(clock), .in1(_331));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7076 (.out1(R7077), .clock(clock), .in1(_320));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7077 (.out1(R7078), .clock(clock), .in1(_349));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7078 (.out1(R7079), .clock(clock), .in1(_329));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7079 (.out1(R7080), .clock(clock), .in1(_318));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7080 (.out1(R7081), .clock(clock), .in1(_311));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7081 (.out1(R7082), .clock(clock), .in1(_377));
  SRAM op363 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_350),.ADR(R7078));
  SRAM op343 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_330),.ADR(R7079));
  SRAM op332 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_319),.ADR(R7080));
  SRAM op325 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_312),.ADR(R7081));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op391 (.out1(_378), .in1(R7068), .in2(R7082));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op392 (.out1(_379), .in1(_378), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op383 (.out1(_370), .in1(R7072), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op372 (.out1(_359), .in1(R7073), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op352 (.out1(_339), .in1(R7075), .in2(64 'd 18446744073709551615));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op326 (.out1(_313), .in1(2 'd 2), .in2(R6650));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op393 (.out1(_380), .in1(_379), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op384 (.out1(_371), .in1(R7069), .in2(_370));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op373 (.out1(_360), .in1(R7070), .in2(_359));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op353 (.out1(_340), .in1(R7071), .in2(_339));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op394 (.out1(_381), .in1(_371), .in2(_380));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op374 (.out1(_361), .in1(_360), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op365 (.out1(_352), .in1(R7074), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op354 (.out1(_341), .in1(_340), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op345 (.out1(_332), .in1(R7076), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op334 (.out1(_321), .in1(R7077), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3737 (.out1(R3738), .clock(clock), .in1(R3737));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3993 (.out1(R3994), .clock(clock), .in1(R3993));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4248 (.out1(R4249), .clock(clock), .in1(R4248));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4493 (.out1(R4494), .clock(clock), .in1(R4493));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4733 (.out1(R4734), .clock(clock), .in1(R4733));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5020 (.out1(R5021), .clock(clock), .in1(R5020));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5252 (.out1(R5253), .clock(clock), .in1(R5252));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5479 (.out1(R5480), .clock(clock), .in1(R5479));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5753 (.out1(R5754), .clock(clock), .in1(R5753));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5971 (.out1(R5972), .clock(clock), .in1(R5971));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6184 (.out1(R6185), .clock(clock), .in1(R6184));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6445 (.out1(R6446), .clock(clock), .in1(R6445));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6650 (.out1(R6651), .clock(clock), .in1(R6650));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6850 (.out1(R6851), .clock(clock), .in1(R6850));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7082 (.out1(R7083), .clock(clock), .in1(_350));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7083 (.out1(R7084), .clock(clock), .in1(_330));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7084 (.out1(R7085), .clock(clock), .in1(_319));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7085 (.out1(R7086), .clock(clock), .in1(_312));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7086 (.out1(R7087), .clock(clock), .in1(_313));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7087 (.out1(R7088), .clock(clock), .in1(_381));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7088 (.out1(R7089), .clock(clock), .in1(_361));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7089 (.out1(R7090), .clock(clock), .in1(_352));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7090 (.out1(R7091), .clock(clock), .in1(_341));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7091 (.out1(R7092), .clock(clock), .in1(_332));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7092 (.out1(R7093), .clock(clock), .in1(_321));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op375 (.out1(_362), .in1(R7089), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op366 (.out1(_353), .in1(R7083), .in2(R7090));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op335 (.out1(_322), .in1(R7085), .in2(R7093));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op395 (.out1(_382), .in1(R7088), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op376 (.out1(_363), .in1(_353), .in2(_362));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op355 (.out1(_342), .in1(R7091), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op346 (.out1(_333), .in1(R7084), .in2(R7092));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op336 (.out1(_323), .in1(_322), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op327 (.out1(_314), .in1(R7087), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op356 (.out1(_343), .in1(_333), .in2(_342));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op396 (.out1(_383), .in1(_382), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op377 (.out1(_364), .in1(_363), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op337 (.out1(_324), .in1(_323), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op328 (.out1(_315), .in1(R7086), .in2(_314));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op397 (.out1(_384), .in1(_364), .in2(_383));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op357 (.out1(_344), .in1(_343), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op338 (.out1(_325), .in1(_315), .in2(_324));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3738 (.out1(R3739), .clock(clock), .in1(R3738));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3994 (.out1(R3995), .clock(clock), .in1(R3994));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4249 (.out1(R4250), .clock(clock), .in1(R4249));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4494 (.out1(R4495), .clock(clock), .in1(R4494));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4734 (.out1(R4735), .clock(clock), .in1(R4734));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5021 (.out1(R5022), .clock(clock), .in1(R5021));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5253 (.out1(R5254), .clock(clock), .in1(R5253));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5480 (.out1(R5481), .clock(clock), .in1(R5480));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5754 (.out1(R5755), .clock(clock), .in1(R5754));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5972 (.out1(R5973), .clock(clock), .in1(R5972));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6185 (.out1(R6186), .clock(clock), .in1(R6185));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6446 (.out1(R6447), .clock(clock), .in1(R6446));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6651 (.out1(R6652), .clock(clock), .in1(R6651));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6851 (.out1(R6852), .clock(clock), .in1(R6851));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7093 (.out1(R7094), .clock(clock), .in1(_384));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7094 (.out1(R7095), .clock(clock), .in1(_344));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7095 (.out1(R7096), .clock(clock), .in1(_325));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op318 (.out1(_305), .in1(R6447));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op358 (.out1(_345), .in1(R7095), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op339 (.out1(_326), .in1(R7096), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op398 (.out1(_385), .in1(R7094), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op359 (.out1(_346), .in1(_326), .in2(_345));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op319 (.out1(_306), .in1(_305), .in2(2 'd 2));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op399 (.out1(_386), .in1(_346), .in2(_385));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op400 (.out1(_387), .in1(_386), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3739 (.out1(R3740), .clock(clock), .in1(R3739));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3995 (.out1(R3996), .clock(clock), .in1(R3995));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4250 (.out1(R4251), .clock(clock), .in1(R4250));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4495 (.out1(R4496), .clock(clock), .in1(R4495));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4735 (.out1(R4736), .clock(clock), .in1(R4735));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5022 (.out1(R5023), .clock(clock), .in1(R5022));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5254 (.out1(R5255), .clock(clock), .in1(R5254));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5481 (.out1(R5482), .clock(clock), .in1(R5481));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5755 (.out1(R5756), .clock(clock), .in1(R5755));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5973 (.out1(R5974), .clock(clock), .in1(R5973));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6186 (.out1(R6187), .clock(clock), .in1(R6186));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6447 (.out1(R6448), .clock(clock), .in1(R6447));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6652 (.out1(R6653), .clock(clock), .in1(R6652));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6852 (.out1(R6853), .clock(clock), .in1(R6852));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7096 (.out1(R7097), .clock(clock), .in1(_306));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7097 (.out1(R7098), .clock(clock), .in1(_387));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op401 (.out1(_388), .in1(R7098), .in2(57 'd 72340172838076673));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op320 (.out1(_307), .in1(base0_34_3568_D), .in2(R7097));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3740 (.out1(R3741), .clock(clock), .in1(R3740));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3996 (.out1(R3997), .clock(clock), .in1(R3996));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4251 (.out1(R4252), .clock(clock), .in1(R4251));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4496 (.out1(R4497), .clock(clock), .in1(R4496));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4736 (.out1(R4737), .clock(clock), .in1(R4736));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5023 (.out1(R5024), .clock(clock), .in1(R5023));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5255 (.out1(R5256), .clock(clock), .in1(R5255));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5482 (.out1(R5483), .clock(clock), .in1(R5482));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5756 (.out1(R5757), .clock(clock), .in1(R5756));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5974 (.out1(R5975), .clock(clock), .in1(R5974));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6187 (.out1(R6188), .clock(clock), .in1(R6187));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6448 (.out1(R6449), .clock(clock), .in1(R6448));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6653 (.out1(R6654), .clock(clock), .in1(R6653));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6853 (.out1(R6854), .clock(clock), .in1(R6853));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7098 (.out1(R7099), .clock(clock), .in1(_388));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7099 (.out1(R7100), .clock(clock), .in1(_307));
  SRAM op321 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_308),.ADR(R7100));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op402 (.out1(_389), .in1(R7099), .in2(6 'd 56));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3741 (.out1(R3742), .clock(clock), .in1(R3741));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3997 (.out1(R3998), .clock(clock), .in1(R3997));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4252 (.out1(R4253), .clock(clock), .in1(R4252));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4497 (.out1(R4498), .clock(clock), .in1(R4497));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4737 (.out1(R4738), .clock(clock), .in1(R4737));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5024 (.out1(R5025), .clock(clock), .in1(R5024));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5256 (.out1(R5257), .clock(clock), .in1(R5256));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5483 (.out1(R5484), .clock(clock), .in1(R5483));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5757 (.out1(R5758), .clock(clock), .in1(R5757));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5975 (.out1(R5976), .clock(clock), .in1(R5975));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6188 (.out1(R6189), .clock(clock), .in1(R6188));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6449 (.out1(R6450), .clock(clock), .in1(R6449));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6654 (.out1(R6655), .clock(clock), .in1(R6654));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6854 (.out1(R6855), .clock(clock), .in1(R6854));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7100 (.out1(R7101), .clock(clock), .in1(_308));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7101 (.out1(R7102), .clock(clock), .in1(_389));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op403 (.out1(_390), .in1(R7102));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op404 (.out1(_391), .in1(R7101), .in2(_390));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op405 (.out1(idx_3569), .in1(_391), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3742 (.out1(R3743), .clock(clock), .in1(R3742));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3998 (.out1(R3999), .clock(clock), .in1(R3998));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4253 (.out1(R4254), .clock(clock), .in1(R4253));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4498 (.out1(R4499), .clock(clock), .in1(R4498));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4738 (.out1(R4739), .clock(clock), .in1(R4738));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5025 (.out1(R5026), .clock(clock), .in1(R5025));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5257 (.out1(R5258), .clock(clock), .in1(R5257));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5484 (.out1(R5485), .clock(clock), .in1(R5484));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5758 (.out1(R5759), .clock(clock), .in1(R5758));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5976 (.out1(R5977), .clock(clock), .in1(R5976));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6189 (.out1(R6190), .clock(clock), .in1(R6189));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6450 (.out1(R6451), .clock(clock), .in1(R6450));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6655 (.out1(R6656), .clock(clock), .in1(R6655));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6855 (.out1(R6856), .clock(clock), .in1(R6855));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7102 (.out1(R7103), .clock(clock), .in1(idx_3569));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op409 (.out1(_394), .in1(R7103));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op410 (.out1(_395), .in1(_394), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3743 (.out1(R3744), .clock(clock), .in1(R3743));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op3999 (.out1(R4000), .clock(clock), .in1(R3999));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4254 (.out1(R4255), .clock(clock), .in1(R4254));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4499 (.out1(R4500), .clock(clock), .in1(R4499));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4739 (.out1(R4740), .clock(clock), .in1(R4739));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5026 (.out1(R5027), .clock(clock), .in1(R5026));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5258 (.out1(R5259), .clock(clock), .in1(R5258));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5485 (.out1(R5486), .clock(clock), .in1(R5485));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5759 (.out1(R5760), .clock(clock), .in1(R5759));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5977 (.out1(R5978), .clock(clock), .in1(R5977));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6190 (.out1(R6191), .clock(clock), .in1(R6190));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6451 (.out1(R6452), .clock(clock), .in1(R6451));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6656 (.out1(R6657), .clock(clock), .in1(R6656));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6856 (.out1(R6857), .clock(clock), .in1(R6856));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7103 (.out1(R7104), .clock(clock), .in1(R7103));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7295 (.out1(R7296), .clock(clock), .in1(_395));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op411 (.out1(_396), .in1(vec40_3571_D), .in2(R7296));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3744 (.out1(R3745), .clock(clock), .in1(R3744));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4000 (.out1(R4001), .clock(clock), .in1(R4000));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4255 (.out1(R4256), .clock(clock), .in1(R4255));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4500 (.out1(R4501), .clock(clock), .in1(R4500));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4740 (.out1(R4741), .clock(clock), .in1(R4740));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5027 (.out1(R5028), .clock(clock), .in1(R5027));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5259 (.out1(R5260), .clock(clock), .in1(R5259));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5486 (.out1(R5487), .clock(clock), .in1(R5486));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5760 (.out1(R5761), .clock(clock), .in1(R5760));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5978 (.out1(R5979), .clock(clock), .in1(R5978));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6191 (.out1(R6192), .clock(clock), .in1(R6191));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6452 (.out1(R6453), .clock(clock), .in1(R6452));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6657 (.out1(R6658), .clock(clock), .in1(R6657));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6857 (.out1(R6858), .clock(clock), .in1(R6857));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7104 (.out1(R7105), .clock(clock), .in1(R7104));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7296 (.out1(R7297), .clock(clock), .in1(_396));
  SRAM op412 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_397),.ADR(R7297));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3745 (.out1(R3746), .clock(clock), .in1(R3745));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4001 (.out1(R4002), .clock(clock), .in1(R4001));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4256 (.out1(R4257), .clock(clock), .in1(R4256));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4501 (.out1(R4502), .clock(clock), .in1(R4501));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4741 (.out1(R4742), .clock(clock), .in1(R4741));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5028 (.out1(R5029), .clock(clock), .in1(R5028));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5260 (.out1(R5261), .clock(clock), .in1(R5260));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5487 (.out1(R5488), .clock(clock), .in1(R5487));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5761 (.out1(R5762), .clock(clock), .in1(R5761));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5979 (.out1(R5980), .clock(clock), .in1(R5979));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6192 (.out1(R6193), .clock(clock), .in1(R6192));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6453 (.out1(R6454), .clock(clock), .in1(R6453));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6658 (.out1(R6659), .clock(clock), .in1(R6658));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6858 (.out1(R6859), .clock(clock), .in1(R6858));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7105 (.out1(R7106), .clock(clock), .in1(R7105));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7297 (.out1(R7298), .clock(clock), .in1(_397));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(5), .BITSIZE_out1(64), .PRECISION(64)) op406 (.out1(_392), .in1(ip1_3530_D), .in2(5 'd 18));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op407 (.out1(_393), .in1(_392));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op408 (.out1(off_3570), .in1(_393), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op413 (.out1(_398), .in1(R7298), .in2(off_3570));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3746 (.out1(R3747), .clock(clock), .in1(R3746));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4002 (.out1(R4003), .clock(clock), .in1(R4002));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4257 (.out1(R4258), .clock(clock), .in1(R4257));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4502 (.out1(R4503), .clock(clock), .in1(R4502));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4742 (.out1(R4743), .clock(clock), .in1(R4742));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5029 (.out1(R5030), .clock(clock), .in1(R5029));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5261 (.out1(R5262), .clock(clock), .in1(R5261));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5488 (.out1(R5489), .clock(clock), .in1(R5488));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5762 (.out1(R5763), .clock(clock), .in1(R5762));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5980 (.out1(R5981), .clock(clock), .in1(R5980));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6193 (.out1(R6194), .clock(clock), .in1(R6193));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6454 (.out1(R6455), .clock(clock), .in1(R6454));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6659 (.out1(R6660), .clock(clock), .in1(R6659));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6859 (.out1(R6860), .clock(clock), .in1(R6859));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7106 (.out1(R7107), .clock(clock), .in1(R7106));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7298 (.out1(R7299), .clock(clock), .in1(off_3570));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7485 (.out1(R7486), .clock(clock), .in1(_398));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op414 (.out1(_399), .in1(R7486), .in2(1 'd 1));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op415 (.out1(ifout415), .in1(_399), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op483 (.out1(_467), .in1(R7107));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op476 (.out1(_460), .in1(R7107));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op465 (.out1(_449), .in1(R7107));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op445 (.out1(_429), .in1(R7107));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op484 (.out1(_468), .in1(_467), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op477 (.out1(_461), .in1(_460), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op466 (.out1(_450), .in1(_449), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op446 (.out1(_430), .in1(_429), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3747 (.out1(R3748), .clock(clock), .in1(R3747));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4003 (.out1(R4004), .clock(clock), .in1(R4003));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4258 (.out1(R4259), .clock(clock), .in1(R4258));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4503 (.out1(R4504), .clock(clock), .in1(R4503));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4743 (.out1(R4744), .clock(clock), .in1(R4743));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5030 (.out1(R5031), .clock(clock), .in1(R5030));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5262 (.out1(R5263), .clock(clock), .in1(R5262));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5489 (.out1(R5490), .clock(clock), .in1(R5489));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5763 (.out1(R5764), .clock(clock), .in1(R5763));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5981 (.out1(R5982), .clock(clock), .in1(R5981));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6194 (.out1(R6195), .clock(clock), .in1(R6194));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6455 (.out1(R6456), .clock(clock), .in1(R6455));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6660 (.out1(R6661), .clock(clock), .in1(R6660));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6860 (.out1(R6861), .clock(clock), .in1(R6860));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7107 (.out1(R7108), .clock(clock), .in1(R7107));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7299 (.out1(R7300), .clock(clock), .in1(R7299));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7486 (.out1(R7487), .clock(clock), .in1(ifout415));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7680 (.out1(R7681), .clock(clock), .in1(_468));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7681 (.out1(R7682), .clock(clock), .in1(_461));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7682 (.out1(R7683), .clock(clock), .in1(_450));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7683 (.out1(R7684), .clock(clock), .in1(_430));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op458 (.out1(_442), .in1(R7108));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op438 (.out1(_422), .in1(R7108));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op427 (.out1(_411), .in1(R7108));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op420 (.out1(_404), .in1(R7108));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op487 (.out1(_471), .in1(2 'd 2), .in2(R7300));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op459 (.out1(_443), .in1(_442), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op439 (.out1(_423), .in1(_422), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op428 (.out1(_412), .in1(_411), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op421 (.out1(_405), .in1(_404), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op485 (.out1(_469), .in1(vec40_3571_D), .in2(R7681));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op478 (.out1(_462), .in1(vec40_3571_D), .in2(R7682));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op467 (.out1(_451), .in1(vec40_3571_D), .in2(R7683));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op447 (.out1(_431), .in1(vec40_3571_D), .in2(R7684));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3748 (.out1(R3749), .clock(clock), .in1(R3748));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4004 (.out1(R4005), .clock(clock), .in1(R4004));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4259 (.out1(R4260), .clock(clock), .in1(R4259));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4504 (.out1(R4505), .clock(clock), .in1(R4504));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4744 (.out1(R4745), .clock(clock), .in1(R4744));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5031 (.out1(R5032), .clock(clock), .in1(R5031));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5263 (.out1(R5264), .clock(clock), .in1(R5263));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5490 (.out1(R5491), .clock(clock), .in1(R5490));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5764 (.out1(R5765), .clock(clock), .in1(R5764));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5982 (.out1(R5983), .clock(clock), .in1(R5982));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6195 (.out1(R6196), .clock(clock), .in1(R6195));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6456 (.out1(R6457), .clock(clock), .in1(R6456));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6661 (.out1(R6662), .clock(clock), .in1(R6661));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6861 (.out1(R6862), .clock(clock), .in1(R6861));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7108 (.out1(R7109), .clock(clock), .in1(R7108));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7300 (.out1(R7301), .clock(clock), .in1(R7300));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7487 (.out1(R7488), .clock(clock), .in1(R7487));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7684 (.out1(R7685), .clock(clock), .in1(_471));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7685 (.out1(R7686), .clock(clock), .in1(_443));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7686 (.out1(R7687), .clock(clock), .in1(_423));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7687 (.out1(R7688), .clock(clock), .in1(_412));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7688 (.out1(R7689), .clock(clock), .in1(_405));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7689 (.out1(R7690), .clock(clock), .in1(_469));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7690 (.out1(R7691), .clock(clock), .in1(_462));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7691 (.out1(R7692), .clock(clock), .in1(_451));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7692 (.out1(R7693), .clock(clock), .in1(_431));
  SRAM op486 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_470),.ADR(R7690));
  SRAM op479 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_463),.ADR(R7691));
  SRAM op468 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_452),.ADR(R7692));
  SRAM op448 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_432),.ADR(R7693));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op480 (.out1(_464), .in1(2 'd 2), .in2(R7301));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op469 (.out1(_453), .in1(2 'd 2), .in2(R7301));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op462 (.out1(_446), .in1(2 'd 2), .in2(R7301));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op449 (.out1(_433), .in1(2 'd 2), .in2(R7301));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op442 (.out1(_426), .in1(2 'd 2), .in2(R7301));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op431 (.out1(_415), .in1(2 'd 2), .in2(R7301));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op460 (.out1(_444), .in1(vec40_3571_D), .in2(R7686));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op440 (.out1(_424), .in1(vec40_3571_D), .in2(R7687));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op429 (.out1(_413), .in1(vec40_3571_D), .in2(R7688));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op422 (.out1(_406), .in1(vec40_3571_D), .in2(R7689));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op488 (.out1(_472), .in1(R7685), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3749 (.out1(R3750), .clock(clock), .in1(R3749));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4005 (.out1(R4006), .clock(clock), .in1(R4005));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4260 (.out1(R4261), .clock(clock), .in1(R4260));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4505 (.out1(R4506), .clock(clock), .in1(R4505));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4745 (.out1(R4746), .clock(clock), .in1(R4745));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5032 (.out1(R5033), .clock(clock), .in1(R5032));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5264 (.out1(R5265), .clock(clock), .in1(R5264));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5491 (.out1(R5492), .clock(clock), .in1(R5491));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5765 (.out1(R5766), .clock(clock), .in1(R5765));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5983 (.out1(R5984), .clock(clock), .in1(R5983));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6196 (.out1(R6197), .clock(clock), .in1(R6196));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6457 (.out1(R6458), .clock(clock), .in1(R6457));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6662 (.out1(R6663), .clock(clock), .in1(R6662));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6862 (.out1(R6863), .clock(clock), .in1(R6862));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7109 (.out1(R7110), .clock(clock), .in1(R7109));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7301 (.out1(R7302), .clock(clock), .in1(R7301));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7488 (.out1(R7489), .clock(clock), .in1(R7488));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7693 (.out1(R7694), .clock(clock), .in1(_470));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7694 (.out1(R7695), .clock(clock), .in1(_463));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7695 (.out1(R7696), .clock(clock), .in1(_452));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7696 (.out1(R7697), .clock(clock), .in1(_432));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7697 (.out1(R7698), .clock(clock), .in1(_464));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7698 (.out1(R7699), .clock(clock), .in1(_453));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7699 (.out1(R7700), .clock(clock), .in1(_446));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7700 (.out1(R7701), .clock(clock), .in1(_433));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7701 (.out1(R7702), .clock(clock), .in1(_426));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7702 (.out1(R7703), .clock(clock), .in1(_415));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7703 (.out1(R7704), .clock(clock), .in1(_444));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7704 (.out1(R7705), .clock(clock), .in1(_424));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7705 (.out1(R7706), .clock(clock), .in1(_413));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7706 (.out1(R7707), .clock(clock), .in1(_406));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7707 (.out1(R7708), .clock(clock), .in1(_472));
  SRAM op461 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_445),.ADR(R7704));
  SRAM op441 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_425),.ADR(R7705));
  SRAM op430 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_414),.ADR(R7706));
  SRAM op423 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_407),.ADR(R7707));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op489 (.out1(_473), .in1(R7694), .in2(R7708));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op490 (.out1(_474), .in1(_473), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op481 (.out1(_465), .in1(R7698), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op470 (.out1(_454), .in1(R7699), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op450 (.out1(_434), .in1(R7701), .in2(64 'd 18446744073709551615));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op424 (.out1(_408), .in1(2 'd 2), .in2(R7302));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op491 (.out1(_475), .in1(_474), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op482 (.out1(_466), .in1(R7695), .in2(_465));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op471 (.out1(_455), .in1(R7696), .in2(_454));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op451 (.out1(_435), .in1(R7697), .in2(_434));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op492 (.out1(_476), .in1(_466), .in2(_475));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op472 (.out1(_456), .in1(_455), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op463 (.out1(_447), .in1(R7700), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op452 (.out1(_436), .in1(_435), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op443 (.out1(_427), .in1(R7702), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op432 (.out1(_416), .in1(R7703), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3750 (.out1(R3751), .clock(clock), .in1(R3750));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4006 (.out1(R4007), .clock(clock), .in1(R4006));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4261 (.out1(R4262), .clock(clock), .in1(R4261));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4506 (.out1(R4507), .clock(clock), .in1(R4506));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4746 (.out1(R4747), .clock(clock), .in1(R4746));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5033 (.out1(R5034), .clock(clock), .in1(R5033));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5265 (.out1(R5266), .clock(clock), .in1(R5265));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5492 (.out1(R5493), .clock(clock), .in1(R5492));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5766 (.out1(R5767), .clock(clock), .in1(R5766));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5984 (.out1(R5985), .clock(clock), .in1(R5984));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6197 (.out1(R6198), .clock(clock), .in1(R6197));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6458 (.out1(R6459), .clock(clock), .in1(R6458));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6663 (.out1(R6664), .clock(clock), .in1(R6663));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6863 (.out1(R6864), .clock(clock), .in1(R6863));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7110 (.out1(R7111), .clock(clock), .in1(R7110));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7302 (.out1(R7303), .clock(clock), .in1(R7302));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7489 (.out1(R7490), .clock(clock), .in1(R7489));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7708 (.out1(R7709), .clock(clock), .in1(_445));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7709 (.out1(R7710), .clock(clock), .in1(_425));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7710 (.out1(R7711), .clock(clock), .in1(_414));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7711 (.out1(R7712), .clock(clock), .in1(_407));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7712 (.out1(R7713), .clock(clock), .in1(_408));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7713 (.out1(R7714), .clock(clock), .in1(_476));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7714 (.out1(R7715), .clock(clock), .in1(_456));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7715 (.out1(R7716), .clock(clock), .in1(_447));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7716 (.out1(R7717), .clock(clock), .in1(_436));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7717 (.out1(R7718), .clock(clock), .in1(_427));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7718 (.out1(R7719), .clock(clock), .in1(_416));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op473 (.out1(_457), .in1(R7715), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op464 (.out1(_448), .in1(R7709), .in2(R7716));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op433 (.out1(_417), .in1(R7711), .in2(R7719));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op493 (.out1(_477), .in1(R7714), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op474 (.out1(_458), .in1(_448), .in2(_457));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op453 (.out1(_437), .in1(R7717), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op444 (.out1(_428), .in1(R7710), .in2(R7718));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op434 (.out1(_418), .in1(_417), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op425 (.out1(_409), .in1(R7713), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op454 (.out1(_438), .in1(_428), .in2(_437));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op494 (.out1(_478), .in1(_477), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op475 (.out1(_459), .in1(_458), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op435 (.out1(_419), .in1(_418), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op426 (.out1(_410), .in1(R7712), .in2(_409));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op495 (.out1(_479), .in1(_459), .in2(_478));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op455 (.out1(_439), .in1(_438), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op436 (.out1(_420), .in1(_410), .in2(_419));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3751 (.out1(R3752), .clock(clock), .in1(R3751));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4007 (.out1(R4008), .clock(clock), .in1(R4007));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4262 (.out1(R4263), .clock(clock), .in1(R4262));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4507 (.out1(R4508), .clock(clock), .in1(R4507));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4747 (.out1(R4748), .clock(clock), .in1(R4747));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5034 (.out1(R5035), .clock(clock), .in1(R5034));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5266 (.out1(R5267), .clock(clock), .in1(R5266));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5493 (.out1(R5494), .clock(clock), .in1(R5493));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5767 (.out1(R5768), .clock(clock), .in1(R5767));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5985 (.out1(R5986), .clock(clock), .in1(R5985));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6198 (.out1(R6199), .clock(clock), .in1(R6198));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6459 (.out1(R6460), .clock(clock), .in1(R6459));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6664 (.out1(R6665), .clock(clock), .in1(R6664));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6864 (.out1(R6865), .clock(clock), .in1(R6864));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7111 (.out1(R7112), .clock(clock), .in1(R7111));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7303 (.out1(R7304), .clock(clock), .in1(R7303));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7490 (.out1(R7491), .clock(clock), .in1(R7490));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7719 (.out1(R7720), .clock(clock), .in1(_479));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7720 (.out1(R7721), .clock(clock), .in1(_439));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7721 (.out1(R7722), .clock(clock), .in1(_420));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op416 (.out1(_400), .in1(R7112));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op456 (.out1(_440), .in1(R7721), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op437 (.out1(_421), .in1(R7722), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op496 (.out1(_480), .in1(R7720), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op457 (.out1(_441), .in1(_421), .in2(_440));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op417 (.out1(_401), .in1(_400), .in2(2 'd 2));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op497 (.out1(_481), .in1(_441), .in2(_480));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op498 (.out1(_482), .in1(_481), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3752 (.out1(R3753), .clock(clock), .in1(R3752));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4008 (.out1(R4009), .clock(clock), .in1(R4008));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4263 (.out1(R4264), .clock(clock), .in1(R4263));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4508 (.out1(R4509), .clock(clock), .in1(R4508));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4748 (.out1(R4749), .clock(clock), .in1(R4748));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5035 (.out1(R5036), .clock(clock), .in1(R5035));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5267 (.out1(R5268), .clock(clock), .in1(R5267));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5494 (.out1(R5495), .clock(clock), .in1(R5494));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5768 (.out1(R5769), .clock(clock), .in1(R5768));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5986 (.out1(R5987), .clock(clock), .in1(R5986));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6199 (.out1(R6200), .clock(clock), .in1(R6199));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6460 (.out1(R6461), .clock(clock), .in1(R6460));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6665 (.out1(R6666), .clock(clock), .in1(R6665));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6865 (.out1(R6866), .clock(clock), .in1(R6865));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7112 (.out1(R7113), .clock(clock), .in1(R7112));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7304 (.out1(R7305), .clock(clock), .in1(R7304));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7491 (.out1(R7492), .clock(clock), .in1(R7491));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7722 (.out1(R7723), .clock(clock), .in1(_401));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7723 (.out1(R7724), .clock(clock), .in1(_482));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op499 (.out1(_483), .in1(R7724), .in2(57 'd 72340172838076673));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op418 (.out1(_402), .in1(base0_40_3576_D), .in2(R7723));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3753 (.out1(R3754), .clock(clock), .in1(R3753));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4009 (.out1(R4010), .clock(clock), .in1(R4009));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4264 (.out1(R4265), .clock(clock), .in1(R4264));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4509 (.out1(R4510), .clock(clock), .in1(R4509));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4749 (.out1(R4750), .clock(clock), .in1(R4749));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5036 (.out1(R5037), .clock(clock), .in1(R5036));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5268 (.out1(R5269), .clock(clock), .in1(R5268));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5495 (.out1(R5496), .clock(clock), .in1(R5495));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5769 (.out1(R5770), .clock(clock), .in1(R5769));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5987 (.out1(R5988), .clock(clock), .in1(R5987));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6200 (.out1(R6201), .clock(clock), .in1(R6200));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6461 (.out1(R6462), .clock(clock), .in1(R6461));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6666 (.out1(R6667), .clock(clock), .in1(R6666));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6866 (.out1(R6867), .clock(clock), .in1(R6866));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7113 (.out1(R7114), .clock(clock), .in1(R7113));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7305 (.out1(R7306), .clock(clock), .in1(R7305));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7492 (.out1(R7493), .clock(clock), .in1(R7492));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7724 (.out1(R7725), .clock(clock), .in1(_483));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7725 (.out1(R7726), .clock(clock), .in1(_402));
  SRAM op419 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_403),.ADR(R7726));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op500 (.out1(_484), .in1(R7725), .in2(6 'd 56));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3754 (.out1(R3755), .clock(clock), .in1(R3754));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4010 (.out1(R4011), .clock(clock), .in1(R4010));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4265 (.out1(R4266), .clock(clock), .in1(R4265));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4510 (.out1(R4511), .clock(clock), .in1(R4510));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4750 (.out1(R4751), .clock(clock), .in1(R4750));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5037 (.out1(R5038), .clock(clock), .in1(R5037));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5269 (.out1(R5270), .clock(clock), .in1(R5269));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5496 (.out1(R5497), .clock(clock), .in1(R5496));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5770 (.out1(R5771), .clock(clock), .in1(R5770));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5988 (.out1(R5989), .clock(clock), .in1(R5988));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6201 (.out1(R6202), .clock(clock), .in1(R6201));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6462 (.out1(R6463), .clock(clock), .in1(R6462));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6667 (.out1(R6668), .clock(clock), .in1(R6667));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6867 (.out1(R6868), .clock(clock), .in1(R6867));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7114 (.out1(R7115), .clock(clock), .in1(R7114));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7306 (.out1(R7307), .clock(clock), .in1(R7306));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7493 (.out1(R7494), .clock(clock), .in1(R7493));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7726 (.out1(R7727), .clock(clock), .in1(_403));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7727 (.out1(R7728), .clock(clock), .in1(_484));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op501 (.out1(_485), .in1(R7728));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op502 (.out1(_486), .in1(R7727), .in2(_485));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op503 (.out1(idx_3577), .in1(_486), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3755 (.out1(R3756), .clock(clock), .in1(R3755));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4011 (.out1(R4012), .clock(clock), .in1(R4011));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4266 (.out1(R4267), .clock(clock), .in1(R4266));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4511 (.out1(R4512), .clock(clock), .in1(R4511));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4751 (.out1(R4752), .clock(clock), .in1(R4751));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5038 (.out1(R5039), .clock(clock), .in1(R5038));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5270 (.out1(R5271), .clock(clock), .in1(R5270));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5497 (.out1(R5498), .clock(clock), .in1(R5497));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5771 (.out1(R5772), .clock(clock), .in1(R5771));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5989 (.out1(R5990), .clock(clock), .in1(R5989));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6202 (.out1(R6203), .clock(clock), .in1(R6202));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6463 (.out1(R6464), .clock(clock), .in1(R6463));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6668 (.out1(R6669), .clock(clock), .in1(R6668));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6868 (.out1(R6869), .clock(clock), .in1(R6868));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7115 (.out1(R7116), .clock(clock), .in1(R7115));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7307 (.out1(R7308), .clock(clock), .in1(R7307));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7494 (.out1(R7495), .clock(clock), .in1(R7494));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7728 (.out1(R7729), .clock(clock), .in1(idx_3577));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op507 (.out1(_489), .in1(R7729));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op508 (.out1(_490), .in1(_489), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3756 (.out1(R3757), .clock(clock), .in1(R3756));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4012 (.out1(R4013), .clock(clock), .in1(R4012));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4267 (.out1(R4268), .clock(clock), .in1(R4267));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4512 (.out1(R4513), .clock(clock), .in1(R4512));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4752 (.out1(R4753), .clock(clock), .in1(R4752));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5039 (.out1(R5040), .clock(clock), .in1(R5039));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5271 (.out1(R5272), .clock(clock), .in1(R5271));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5498 (.out1(R5499), .clock(clock), .in1(R5498));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5772 (.out1(R5773), .clock(clock), .in1(R5772));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5990 (.out1(R5991), .clock(clock), .in1(R5990));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6203 (.out1(R6204), .clock(clock), .in1(R6203));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6464 (.out1(R6465), .clock(clock), .in1(R6464));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6669 (.out1(R6670), .clock(clock), .in1(R6669));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6869 (.out1(R6870), .clock(clock), .in1(R6869));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7116 (.out1(R7117), .clock(clock), .in1(R7116));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7308 (.out1(R7309), .clock(clock), .in1(R7308));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7495 (.out1(R7496), .clock(clock), .in1(R7495));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7729 (.out1(R7730), .clock(clock), .in1(R7729));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7908 (.out1(R7909), .clock(clock), .in1(_490));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op509 (.out1(_491), .in1(vec46_3579_D), .in2(R7909));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3757 (.out1(R3758), .clock(clock), .in1(R3757));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4013 (.out1(R4014), .clock(clock), .in1(R4013));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4268 (.out1(R4269), .clock(clock), .in1(R4268));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4513 (.out1(R4514), .clock(clock), .in1(R4513));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4753 (.out1(R4754), .clock(clock), .in1(R4753));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5040 (.out1(R5041), .clock(clock), .in1(R5040));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5272 (.out1(R5273), .clock(clock), .in1(R5272));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5499 (.out1(R5500), .clock(clock), .in1(R5499));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5773 (.out1(R5774), .clock(clock), .in1(R5773));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5991 (.out1(R5992), .clock(clock), .in1(R5991));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6204 (.out1(R6205), .clock(clock), .in1(R6204));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6465 (.out1(R6466), .clock(clock), .in1(R6465));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6670 (.out1(R6671), .clock(clock), .in1(R6670));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6870 (.out1(R6871), .clock(clock), .in1(R6870));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7117 (.out1(R7118), .clock(clock), .in1(R7117));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7309 (.out1(R7310), .clock(clock), .in1(R7309));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7496 (.out1(R7497), .clock(clock), .in1(R7496));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7730 (.out1(R7731), .clock(clock), .in1(R7730));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7909 (.out1(R7910), .clock(clock), .in1(_491));
  SRAM op510 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_492),.ADR(R7910));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3758 (.out1(R3759), .clock(clock), .in1(R3758));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4014 (.out1(R4015), .clock(clock), .in1(R4014));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4269 (.out1(R4270), .clock(clock), .in1(R4269));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4514 (.out1(R4515), .clock(clock), .in1(R4514));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4754 (.out1(R4755), .clock(clock), .in1(R4754));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5041 (.out1(R5042), .clock(clock), .in1(R5041));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5273 (.out1(R5274), .clock(clock), .in1(R5273));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5500 (.out1(R5501), .clock(clock), .in1(R5500));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5774 (.out1(R5775), .clock(clock), .in1(R5774));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5992 (.out1(R5993), .clock(clock), .in1(R5992));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6205 (.out1(R6206), .clock(clock), .in1(R6205));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6466 (.out1(R6467), .clock(clock), .in1(R6466));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6671 (.out1(R6672), .clock(clock), .in1(R6671));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6871 (.out1(R6872), .clock(clock), .in1(R6871));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7118 (.out1(R7119), .clock(clock), .in1(R7118));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7310 (.out1(R7311), .clock(clock), .in1(R7310));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7497 (.out1(R7498), .clock(clock), .in1(R7497));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7731 (.out1(R7732), .clock(clock), .in1(R7731));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op7910 (.out1(R7911), .clock(clock), .in1(_492));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(4), .BITSIZE_out1(64), .PRECISION(64)) op504 (.out1(_487), .in1(ip1_3530_D), .in2(4 'd 12));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op505 (.out1(_488), .in1(_487));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op506 (.out1(off_3578), .in1(_488), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op511 (.out1(_493), .in1(R7911), .in2(off_3578));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3759 (.out1(R3760), .clock(clock), .in1(R3759));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4015 (.out1(R4016), .clock(clock), .in1(R4015));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4270 (.out1(R4271), .clock(clock), .in1(R4270));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4515 (.out1(R4516), .clock(clock), .in1(R4515));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4755 (.out1(R4756), .clock(clock), .in1(R4755));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5042 (.out1(R5043), .clock(clock), .in1(R5042));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5274 (.out1(R5275), .clock(clock), .in1(R5274));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5501 (.out1(R5502), .clock(clock), .in1(R5501));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5775 (.out1(R5776), .clock(clock), .in1(R5775));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5993 (.out1(R5994), .clock(clock), .in1(R5993));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6206 (.out1(R6207), .clock(clock), .in1(R6206));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6467 (.out1(R6468), .clock(clock), .in1(R6467));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6672 (.out1(R6673), .clock(clock), .in1(R6672));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6872 (.out1(R6873), .clock(clock), .in1(R6872));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7119 (.out1(R7120), .clock(clock), .in1(R7119));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7311 (.out1(R7312), .clock(clock), .in1(R7311));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7498 (.out1(R7499), .clock(clock), .in1(R7498));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7732 (.out1(R7733), .clock(clock), .in1(R7732));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7911 (.out1(R7912), .clock(clock), .in1(off_3578));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8085 (.out1(R8086), .clock(clock), .in1(_493));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op512 (.out1(_494), .in1(R8086), .in2(1 'd 1));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op513 (.out1(ifout513), .in1(_494), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op581 (.out1(_562), .in1(R7733));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op574 (.out1(_555), .in1(R7733));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op563 (.out1(_544), .in1(R7733));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op543 (.out1(_524), .in1(R7733));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op582 (.out1(_563), .in1(_562), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op575 (.out1(_556), .in1(_555), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op564 (.out1(_545), .in1(_544), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op544 (.out1(_525), .in1(_524), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3760 (.out1(R3761), .clock(clock), .in1(R3760));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4016 (.out1(R4017), .clock(clock), .in1(R4016));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4271 (.out1(R4272), .clock(clock), .in1(R4271));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4516 (.out1(R4517), .clock(clock), .in1(R4516));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4756 (.out1(R4757), .clock(clock), .in1(R4756));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5043 (.out1(R5044), .clock(clock), .in1(R5043));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5275 (.out1(R5276), .clock(clock), .in1(R5275));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5502 (.out1(R5503), .clock(clock), .in1(R5502));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5776 (.out1(R5777), .clock(clock), .in1(R5776));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5994 (.out1(R5995), .clock(clock), .in1(R5994));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6207 (.out1(R6208), .clock(clock), .in1(R6207));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6468 (.out1(R6469), .clock(clock), .in1(R6468));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6673 (.out1(R6674), .clock(clock), .in1(R6673));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6873 (.out1(R6874), .clock(clock), .in1(R6873));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7120 (.out1(R7121), .clock(clock), .in1(R7120));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7312 (.out1(R7313), .clock(clock), .in1(R7312));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7499 (.out1(R7500), .clock(clock), .in1(R7499));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7733 (.out1(R7734), .clock(clock), .in1(R7733));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7912 (.out1(R7913), .clock(clock), .in1(R7912));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8086 (.out1(R8087), .clock(clock), .in1(ifout513));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8267 (.out1(R8268), .clock(clock), .in1(_563));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8268 (.out1(R8269), .clock(clock), .in1(_556));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8269 (.out1(R8270), .clock(clock), .in1(_545));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8270 (.out1(R8271), .clock(clock), .in1(_525));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op556 (.out1(_537), .in1(R7734));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op536 (.out1(_517), .in1(R7734));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op525 (.out1(_506), .in1(R7734));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op518 (.out1(_499), .in1(R7734));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op585 (.out1(_566), .in1(2 'd 2), .in2(R7913));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op557 (.out1(_538), .in1(_537), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op537 (.out1(_518), .in1(_517), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op526 (.out1(_507), .in1(_506), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op519 (.out1(_500), .in1(_499), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op583 (.out1(_564), .in1(vec46_3579_D), .in2(R8268));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op576 (.out1(_557), .in1(vec46_3579_D), .in2(R8269));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op565 (.out1(_546), .in1(vec46_3579_D), .in2(R8270));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op545 (.out1(_526), .in1(vec46_3579_D), .in2(R8271));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3761 (.out1(R3762), .clock(clock), .in1(R3761));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4017 (.out1(R4018), .clock(clock), .in1(R4017));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4272 (.out1(R4273), .clock(clock), .in1(R4272));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4517 (.out1(R4518), .clock(clock), .in1(R4517));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4757 (.out1(R4758), .clock(clock), .in1(R4757));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5044 (.out1(R5045), .clock(clock), .in1(R5044));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5276 (.out1(R5277), .clock(clock), .in1(R5276));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5503 (.out1(R5504), .clock(clock), .in1(R5503));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5777 (.out1(R5778), .clock(clock), .in1(R5777));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5995 (.out1(R5996), .clock(clock), .in1(R5995));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6208 (.out1(R6209), .clock(clock), .in1(R6208));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6469 (.out1(R6470), .clock(clock), .in1(R6469));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6674 (.out1(R6675), .clock(clock), .in1(R6674));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6874 (.out1(R6875), .clock(clock), .in1(R6874));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7121 (.out1(R7122), .clock(clock), .in1(R7121));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7313 (.out1(R7314), .clock(clock), .in1(R7313));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7500 (.out1(R7501), .clock(clock), .in1(R7500));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7734 (.out1(R7735), .clock(clock), .in1(R7734));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7913 (.out1(R7914), .clock(clock), .in1(R7913));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8087 (.out1(R8088), .clock(clock), .in1(R8087));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8271 (.out1(R8272), .clock(clock), .in1(_566));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8272 (.out1(R8273), .clock(clock), .in1(_538));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8273 (.out1(R8274), .clock(clock), .in1(_518));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8274 (.out1(R8275), .clock(clock), .in1(_507));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8275 (.out1(R8276), .clock(clock), .in1(_500));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8276 (.out1(R8277), .clock(clock), .in1(_564));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8277 (.out1(R8278), .clock(clock), .in1(_557));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8278 (.out1(R8279), .clock(clock), .in1(_546));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8279 (.out1(R8280), .clock(clock), .in1(_526));
  SRAM op584 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_565),.ADR(R8277));
  SRAM op577 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_558),.ADR(R8278));
  SRAM op566 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_547),.ADR(R8279));
  SRAM op546 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_527),.ADR(R8280));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op578 (.out1(_559), .in1(2 'd 2), .in2(R7914));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op567 (.out1(_548), .in1(2 'd 2), .in2(R7914));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op560 (.out1(_541), .in1(2 'd 2), .in2(R7914));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op547 (.out1(_528), .in1(2 'd 2), .in2(R7914));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op540 (.out1(_521), .in1(2 'd 2), .in2(R7914));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op529 (.out1(_510), .in1(2 'd 2), .in2(R7914));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op558 (.out1(_539), .in1(vec46_3579_D), .in2(R8273));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op538 (.out1(_519), .in1(vec46_3579_D), .in2(R8274));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op527 (.out1(_508), .in1(vec46_3579_D), .in2(R8275));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op520 (.out1(_501), .in1(vec46_3579_D), .in2(R8276));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op586 (.out1(_567), .in1(R8272), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3762 (.out1(R3763), .clock(clock), .in1(R3762));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4018 (.out1(R4019), .clock(clock), .in1(R4018));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4273 (.out1(R4274), .clock(clock), .in1(R4273));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4518 (.out1(R4519), .clock(clock), .in1(R4518));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4758 (.out1(R4759), .clock(clock), .in1(R4758));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5045 (.out1(R5046), .clock(clock), .in1(R5045));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5277 (.out1(R5278), .clock(clock), .in1(R5277));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5504 (.out1(R5505), .clock(clock), .in1(R5504));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5778 (.out1(R5779), .clock(clock), .in1(R5778));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5996 (.out1(R5997), .clock(clock), .in1(R5996));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6209 (.out1(R6210), .clock(clock), .in1(R6209));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6470 (.out1(R6471), .clock(clock), .in1(R6470));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6675 (.out1(R6676), .clock(clock), .in1(R6675));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6875 (.out1(R6876), .clock(clock), .in1(R6875));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7122 (.out1(R7123), .clock(clock), .in1(R7122));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7314 (.out1(R7315), .clock(clock), .in1(R7314));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7501 (.out1(R7502), .clock(clock), .in1(R7501));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7735 (.out1(R7736), .clock(clock), .in1(R7735));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7914 (.out1(R7915), .clock(clock), .in1(R7914));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8088 (.out1(R8089), .clock(clock), .in1(R8088));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8280 (.out1(R8281), .clock(clock), .in1(_565));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8281 (.out1(R8282), .clock(clock), .in1(_558));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8282 (.out1(R8283), .clock(clock), .in1(_547));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8283 (.out1(R8284), .clock(clock), .in1(_527));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8284 (.out1(R8285), .clock(clock), .in1(_559));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8285 (.out1(R8286), .clock(clock), .in1(_548));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8286 (.out1(R8287), .clock(clock), .in1(_541));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8287 (.out1(R8288), .clock(clock), .in1(_528));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8288 (.out1(R8289), .clock(clock), .in1(_521));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8289 (.out1(R8290), .clock(clock), .in1(_510));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8290 (.out1(R8291), .clock(clock), .in1(_539));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8291 (.out1(R8292), .clock(clock), .in1(_519));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8292 (.out1(R8293), .clock(clock), .in1(_508));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8293 (.out1(R8294), .clock(clock), .in1(_501));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8294 (.out1(R8295), .clock(clock), .in1(_567));
  SRAM op559 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_540),.ADR(R8291));
  SRAM op539 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_520),.ADR(R8292));
  SRAM op528 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_509),.ADR(R8293));
  SRAM op521 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_502),.ADR(R8294));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op587 (.out1(_568), .in1(R8281), .in2(R8295));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op588 (.out1(_569), .in1(_568), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op579 (.out1(_560), .in1(R8285), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op568 (.out1(_549), .in1(R8286), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op548 (.out1(_529), .in1(R8288), .in2(64 'd 18446744073709551615));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op522 (.out1(_503), .in1(2 'd 2), .in2(R7915));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op589 (.out1(_570), .in1(_569), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op580 (.out1(_561), .in1(R8282), .in2(_560));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op569 (.out1(_550), .in1(R8283), .in2(_549));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op549 (.out1(_530), .in1(R8284), .in2(_529));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op590 (.out1(_571), .in1(_561), .in2(_570));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op570 (.out1(_551), .in1(_550), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op561 (.out1(_542), .in1(R8287), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op550 (.out1(_531), .in1(_530), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op541 (.out1(_522), .in1(R8289), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op530 (.out1(_511), .in1(R8290), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3763 (.out1(R3764), .clock(clock), .in1(R3763));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4019 (.out1(R4020), .clock(clock), .in1(R4019));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4274 (.out1(R4275), .clock(clock), .in1(R4274));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4519 (.out1(R4520), .clock(clock), .in1(R4519));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4759 (.out1(R4760), .clock(clock), .in1(R4759));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5046 (.out1(R5047), .clock(clock), .in1(R5046));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5278 (.out1(R5279), .clock(clock), .in1(R5278));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5505 (.out1(R5506), .clock(clock), .in1(R5505));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5779 (.out1(R5780), .clock(clock), .in1(R5779));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5997 (.out1(R5998), .clock(clock), .in1(R5997));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6210 (.out1(R6211), .clock(clock), .in1(R6210));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6471 (.out1(R6472), .clock(clock), .in1(R6471));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6676 (.out1(R6677), .clock(clock), .in1(R6676));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6876 (.out1(R6877), .clock(clock), .in1(R6876));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7123 (.out1(R7124), .clock(clock), .in1(R7123));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7315 (.out1(R7316), .clock(clock), .in1(R7315));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7502 (.out1(R7503), .clock(clock), .in1(R7502));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7736 (.out1(R7737), .clock(clock), .in1(R7736));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7915 (.out1(R7916), .clock(clock), .in1(R7915));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8089 (.out1(R8090), .clock(clock), .in1(R8089));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8295 (.out1(R8296), .clock(clock), .in1(_540));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8296 (.out1(R8297), .clock(clock), .in1(_520));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8297 (.out1(R8298), .clock(clock), .in1(_509));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8298 (.out1(R8299), .clock(clock), .in1(_502));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8299 (.out1(R8300), .clock(clock), .in1(_503));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8300 (.out1(R8301), .clock(clock), .in1(_571));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8301 (.out1(R8302), .clock(clock), .in1(_551));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8302 (.out1(R8303), .clock(clock), .in1(_542));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8303 (.out1(R8304), .clock(clock), .in1(_531));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8304 (.out1(R8305), .clock(clock), .in1(_522));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8305 (.out1(R8306), .clock(clock), .in1(_511));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op571 (.out1(_552), .in1(R8302), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op562 (.out1(_543), .in1(R8296), .in2(R8303));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op531 (.out1(_512), .in1(R8298), .in2(R8306));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op591 (.out1(_572), .in1(R8301), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op572 (.out1(_553), .in1(_543), .in2(_552));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op551 (.out1(_532), .in1(R8304), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op542 (.out1(_523), .in1(R8297), .in2(R8305));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op532 (.out1(_513), .in1(_512), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op523 (.out1(_504), .in1(R8300), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op552 (.out1(_533), .in1(_523), .in2(_532));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op592 (.out1(_573), .in1(_572), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op573 (.out1(_554), .in1(_553), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op533 (.out1(_514), .in1(_513), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op524 (.out1(_505), .in1(R8299), .in2(_504));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op593 (.out1(_574), .in1(_554), .in2(_573));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op553 (.out1(_534), .in1(_533), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op534 (.out1(_515), .in1(_505), .in2(_514));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3764 (.out1(R3765), .clock(clock), .in1(R3764));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4020 (.out1(R4021), .clock(clock), .in1(R4020));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4275 (.out1(R4276), .clock(clock), .in1(R4275));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4520 (.out1(R4521), .clock(clock), .in1(R4520));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4760 (.out1(R4761), .clock(clock), .in1(R4760));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5047 (.out1(R5048), .clock(clock), .in1(R5047));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5279 (.out1(R5280), .clock(clock), .in1(R5279));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5506 (.out1(R5507), .clock(clock), .in1(R5506));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5780 (.out1(R5781), .clock(clock), .in1(R5780));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5998 (.out1(R5999), .clock(clock), .in1(R5998));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6211 (.out1(R6212), .clock(clock), .in1(R6211));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6472 (.out1(R6473), .clock(clock), .in1(R6472));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6677 (.out1(R6678), .clock(clock), .in1(R6677));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6877 (.out1(R6878), .clock(clock), .in1(R6877));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7124 (.out1(R7125), .clock(clock), .in1(R7124));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7316 (.out1(R7317), .clock(clock), .in1(R7316));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7503 (.out1(R7504), .clock(clock), .in1(R7503));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7737 (.out1(R7738), .clock(clock), .in1(R7737));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7916 (.out1(R7917), .clock(clock), .in1(R7916));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8090 (.out1(R8091), .clock(clock), .in1(R8090));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8306 (.out1(R8307), .clock(clock), .in1(_574));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8307 (.out1(R8308), .clock(clock), .in1(_534));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8308 (.out1(R8309), .clock(clock), .in1(_515));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op514 (.out1(_495), .in1(R7738));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op554 (.out1(_535), .in1(R8308), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op535 (.out1(_516), .in1(R8309), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op594 (.out1(_575), .in1(R8307), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op555 (.out1(_536), .in1(_516), .in2(_535));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op515 (.out1(_496), .in1(_495), .in2(2 'd 2));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op595 (.out1(_576), .in1(_536), .in2(_575));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op596 (.out1(_577), .in1(_576), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3765 (.out1(R3766), .clock(clock), .in1(R3765));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4021 (.out1(R4022), .clock(clock), .in1(R4021));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4276 (.out1(R4277), .clock(clock), .in1(R4276));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4521 (.out1(R4522), .clock(clock), .in1(R4521));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4761 (.out1(R4762), .clock(clock), .in1(R4761));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5048 (.out1(R5049), .clock(clock), .in1(R5048));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5280 (.out1(R5281), .clock(clock), .in1(R5280));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5507 (.out1(R5508), .clock(clock), .in1(R5507));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5781 (.out1(R5782), .clock(clock), .in1(R5781));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5999 (.out1(R6000), .clock(clock), .in1(R5999));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6212 (.out1(R6213), .clock(clock), .in1(R6212));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6473 (.out1(R6474), .clock(clock), .in1(R6473));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6678 (.out1(R6679), .clock(clock), .in1(R6678));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6878 (.out1(R6879), .clock(clock), .in1(R6878));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7125 (.out1(R7126), .clock(clock), .in1(R7125));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7317 (.out1(R7318), .clock(clock), .in1(R7317));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7504 (.out1(R7505), .clock(clock), .in1(R7504));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7738 (.out1(R7739), .clock(clock), .in1(R7738));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7917 (.out1(R7918), .clock(clock), .in1(R7917));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8091 (.out1(R8092), .clock(clock), .in1(R8091));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8309 (.out1(R8310), .clock(clock), .in1(_496));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8310 (.out1(R8311), .clock(clock), .in1(_577));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op597 (.out1(_578), .in1(R8311), .in2(57 'd 72340172838076673));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op516 (.out1(_497), .in1(base0_46_3584_D), .in2(R8310));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3766 (.out1(R3767), .clock(clock), .in1(R3766));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4022 (.out1(R4023), .clock(clock), .in1(R4022));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4277 (.out1(R4278), .clock(clock), .in1(R4277));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4522 (.out1(R4523), .clock(clock), .in1(R4522));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4762 (.out1(R4763), .clock(clock), .in1(R4762));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5049 (.out1(R5050), .clock(clock), .in1(R5049));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5281 (.out1(R5282), .clock(clock), .in1(R5281));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5508 (.out1(R5509), .clock(clock), .in1(R5508));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5782 (.out1(R5783), .clock(clock), .in1(R5782));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6000 (.out1(R6001), .clock(clock), .in1(R6000));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6213 (.out1(R6214), .clock(clock), .in1(R6213));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6474 (.out1(R6475), .clock(clock), .in1(R6474));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6679 (.out1(R6680), .clock(clock), .in1(R6679));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6879 (.out1(R6880), .clock(clock), .in1(R6879));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7126 (.out1(R7127), .clock(clock), .in1(R7126));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7318 (.out1(R7319), .clock(clock), .in1(R7318));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7505 (.out1(R7506), .clock(clock), .in1(R7505));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7739 (.out1(R7740), .clock(clock), .in1(R7739));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7918 (.out1(R7919), .clock(clock), .in1(R7918));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8092 (.out1(R8093), .clock(clock), .in1(R8092));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8311 (.out1(R8312), .clock(clock), .in1(_578));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8312 (.out1(R8313), .clock(clock), .in1(_497));
  SRAM op517 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_498),.ADR(R8313));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op598 (.out1(_579), .in1(R8312), .in2(6 'd 56));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3767 (.out1(R3768), .clock(clock), .in1(R3767));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4023 (.out1(R4024), .clock(clock), .in1(R4023));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4278 (.out1(R4279), .clock(clock), .in1(R4278));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4523 (.out1(R4524), .clock(clock), .in1(R4523));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4763 (.out1(R4764), .clock(clock), .in1(R4763));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5050 (.out1(R5051), .clock(clock), .in1(R5050));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5282 (.out1(R5283), .clock(clock), .in1(R5282));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5509 (.out1(R5510), .clock(clock), .in1(R5509));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5783 (.out1(R5784), .clock(clock), .in1(R5783));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6001 (.out1(R6002), .clock(clock), .in1(R6001));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6214 (.out1(R6215), .clock(clock), .in1(R6214));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6475 (.out1(R6476), .clock(clock), .in1(R6475));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6680 (.out1(R6681), .clock(clock), .in1(R6680));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6880 (.out1(R6881), .clock(clock), .in1(R6880));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7127 (.out1(R7128), .clock(clock), .in1(R7127));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7319 (.out1(R7320), .clock(clock), .in1(R7319));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7506 (.out1(R7507), .clock(clock), .in1(R7506));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7740 (.out1(R7741), .clock(clock), .in1(R7740));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7919 (.out1(R7920), .clock(clock), .in1(R7919));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8093 (.out1(R8094), .clock(clock), .in1(R8093));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8313 (.out1(R8314), .clock(clock), .in1(_498));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8314 (.out1(R8315), .clock(clock), .in1(_579));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op599 (.out1(_580), .in1(R8315));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op600 (.out1(_581), .in1(R8314), .in2(_580));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op601 (.out1(idx_3585), .in1(_581), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3768 (.out1(R3769), .clock(clock), .in1(R3768));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4024 (.out1(R4025), .clock(clock), .in1(R4024));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4279 (.out1(R4280), .clock(clock), .in1(R4279));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4524 (.out1(R4525), .clock(clock), .in1(R4524));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4764 (.out1(R4765), .clock(clock), .in1(R4764));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5051 (.out1(R5052), .clock(clock), .in1(R5051));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5283 (.out1(R5284), .clock(clock), .in1(R5283));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5510 (.out1(R5511), .clock(clock), .in1(R5510));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5784 (.out1(R5785), .clock(clock), .in1(R5784));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6002 (.out1(R6003), .clock(clock), .in1(R6002));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6215 (.out1(R6216), .clock(clock), .in1(R6215));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6476 (.out1(R6477), .clock(clock), .in1(R6476));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6681 (.out1(R6682), .clock(clock), .in1(R6681));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6881 (.out1(R6882), .clock(clock), .in1(R6881));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7128 (.out1(R7129), .clock(clock), .in1(R7128));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7320 (.out1(R7321), .clock(clock), .in1(R7320));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7507 (.out1(R7508), .clock(clock), .in1(R7507));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7741 (.out1(R7742), .clock(clock), .in1(R7741));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7920 (.out1(R7921), .clock(clock), .in1(R7920));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8094 (.out1(R8095), .clock(clock), .in1(R8094));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8315 (.out1(R8316), .clock(clock), .in1(idx_3585));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op605 (.out1(_584), .in1(R8316));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op606 (.out1(_585), .in1(_584), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3769 (.out1(R3770), .clock(clock), .in1(R3769));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4025 (.out1(R4026), .clock(clock), .in1(R4025));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4280 (.out1(R4281), .clock(clock), .in1(R4280));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4525 (.out1(R4526), .clock(clock), .in1(R4525));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4765 (.out1(R4766), .clock(clock), .in1(R4765));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5052 (.out1(R5053), .clock(clock), .in1(R5052));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5284 (.out1(R5285), .clock(clock), .in1(R5284));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5511 (.out1(R5512), .clock(clock), .in1(R5511));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5785 (.out1(R5786), .clock(clock), .in1(R5785));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6003 (.out1(R6004), .clock(clock), .in1(R6003));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6216 (.out1(R6217), .clock(clock), .in1(R6216));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6477 (.out1(R6478), .clock(clock), .in1(R6477));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6682 (.out1(R6683), .clock(clock), .in1(R6682));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6882 (.out1(R6883), .clock(clock), .in1(R6882));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7129 (.out1(R7130), .clock(clock), .in1(R7129));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7321 (.out1(R7322), .clock(clock), .in1(R7321));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7508 (.out1(R7509), .clock(clock), .in1(R7508));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7742 (.out1(R7743), .clock(clock), .in1(R7742));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7921 (.out1(R7922), .clock(clock), .in1(R7921));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8095 (.out1(R8096), .clock(clock), .in1(R8095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8316 (.out1(R8317), .clock(clock), .in1(R8316));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8482 (.out1(R8483), .clock(clock), .in1(_585));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op607 (.out1(_586), .in1(vec52_3587_D), .in2(R8483));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3770 (.out1(R3771), .clock(clock), .in1(R3770));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4026 (.out1(R4027), .clock(clock), .in1(R4026));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4281 (.out1(R4282), .clock(clock), .in1(R4281));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4526 (.out1(R4527), .clock(clock), .in1(R4526));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4766 (.out1(R4767), .clock(clock), .in1(R4766));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5053 (.out1(R5054), .clock(clock), .in1(R5053));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5285 (.out1(R5286), .clock(clock), .in1(R5285));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5512 (.out1(R5513), .clock(clock), .in1(R5512));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5786 (.out1(R5787), .clock(clock), .in1(R5786));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6004 (.out1(R6005), .clock(clock), .in1(R6004));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6217 (.out1(R6218), .clock(clock), .in1(R6217));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6478 (.out1(R6479), .clock(clock), .in1(R6478));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6683 (.out1(R6684), .clock(clock), .in1(R6683));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6883 (.out1(R6884), .clock(clock), .in1(R6883));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7130 (.out1(R7131), .clock(clock), .in1(R7130));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7322 (.out1(R7323), .clock(clock), .in1(R7322));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7509 (.out1(R7510), .clock(clock), .in1(R7509));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7743 (.out1(R7744), .clock(clock), .in1(R7743));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7922 (.out1(R7923), .clock(clock), .in1(R7922));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8096 (.out1(R8097), .clock(clock), .in1(R8096));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8317 (.out1(R8318), .clock(clock), .in1(R8317));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8483 (.out1(R8484), .clock(clock), .in1(_586));
  SRAM op608 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_587),.ADR(R8484));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3771 (.out1(R3772), .clock(clock), .in1(R3771));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4027 (.out1(R4028), .clock(clock), .in1(R4027));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4282 (.out1(R4283), .clock(clock), .in1(R4282));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4527 (.out1(R4528), .clock(clock), .in1(R4527));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4767 (.out1(R4768), .clock(clock), .in1(R4767));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5054 (.out1(R5055), .clock(clock), .in1(R5054));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5286 (.out1(R5287), .clock(clock), .in1(R5286));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5513 (.out1(R5514), .clock(clock), .in1(R5513));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5787 (.out1(R5788), .clock(clock), .in1(R5787));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6005 (.out1(R6006), .clock(clock), .in1(R6005));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6218 (.out1(R6219), .clock(clock), .in1(R6218));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6479 (.out1(R6480), .clock(clock), .in1(R6479));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6684 (.out1(R6685), .clock(clock), .in1(R6684));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6884 (.out1(R6885), .clock(clock), .in1(R6884));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7131 (.out1(R7132), .clock(clock), .in1(R7131));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7323 (.out1(R7324), .clock(clock), .in1(R7323));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7510 (.out1(R7511), .clock(clock), .in1(R7510));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7744 (.out1(R7745), .clock(clock), .in1(R7744));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7923 (.out1(R7924), .clock(clock), .in1(R7923));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8097 (.out1(R8098), .clock(clock), .in1(R8097));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8318 (.out1(R8319), .clock(clock), .in1(R8318));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8484 (.out1(R8485), .clock(clock), .in1(_587));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op602 (.out1(_582), .in1(ip1_3530_D), .in2(3 'd 6));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op603 (.out1(_583), .in1(_582));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op604 (.out1(off_3586), .in1(_583), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op609 (.out1(_588), .in1(R8485), .in2(off_3586));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3772 (.out1(R3773), .clock(clock), .in1(R3772));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4028 (.out1(R4029), .clock(clock), .in1(R4028));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4283 (.out1(R4284), .clock(clock), .in1(R4283));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4528 (.out1(R4529), .clock(clock), .in1(R4528));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4768 (.out1(R4769), .clock(clock), .in1(R4768));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5055 (.out1(R5056), .clock(clock), .in1(R5055));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5287 (.out1(R5288), .clock(clock), .in1(R5287));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5514 (.out1(R5515), .clock(clock), .in1(R5514));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5788 (.out1(R5789), .clock(clock), .in1(R5788));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6006 (.out1(R6007), .clock(clock), .in1(R6006));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6219 (.out1(R6220), .clock(clock), .in1(R6219));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6480 (.out1(R6481), .clock(clock), .in1(R6480));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6685 (.out1(R6686), .clock(clock), .in1(R6685));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6885 (.out1(R6886), .clock(clock), .in1(R6885));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7132 (.out1(R7133), .clock(clock), .in1(R7132));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7324 (.out1(R7325), .clock(clock), .in1(R7324));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7511 (.out1(R7512), .clock(clock), .in1(R7511));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7745 (.out1(R7746), .clock(clock), .in1(R7745));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7924 (.out1(R7925), .clock(clock), .in1(R7924));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8098 (.out1(R8099), .clock(clock), .in1(R8098));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8319 (.out1(R8320), .clock(clock), .in1(R8319));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8485 (.out1(R8486), .clock(clock), .in1(off_3586));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8646 (.out1(R8647), .clock(clock), .in1(_588));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op610 (.out1(_589), .in1(R8647), .in2(1 'd 1));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op611 (.out1(ifout611), .in1(_589), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op679 (.out1(_657), .in1(R8320));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op672 (.out1(_650), .in1(R8320));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op661 (.out1(_639), .in1(R8320));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op641 (.out1(_619), .in1(R8320));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op680 (.out1(_658), .in1(_657), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op673 (.out1(_651), .in1(_650), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op662 (.out1(_640), .in1(_639), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op642 (.out1(_620), .in1(_619), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3773 (.out1(R3774), .clock(clock), .in1(R3773));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4029 (.out1(R4030), .clock(clock), .in1(R4029));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4284 (.out1(R4285), .clock(clock), .in1(R4284));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4529 (.out1(R4530), .clock(clock), .in1(R4529));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4769 (.out1(R4770), .clock(clock), .in1(R4769));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5056 (.out1(R5057), .clock(clock), .in1(R5056));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5288 (.out1(R5289), .clock(clock), .in1(R5288));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5515 (.out1(R5516), .clock(clock), .in1(R5515));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5789 (.out1(R5790), .clock(clock), .in1(R5789));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6007 (.out1(R6008), .clock(clock), .in1(R6007));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6220 (.out1(R6221), .clock(clock), .in1(R6220));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6481 (.out1(R6482), .clock(clock), .in1(R6481));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6686 (.out1(R6687), .clock(clock), .in1(R6686));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6886 (.out1(R6887), .clock(clock), .in1(R6886));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7133 (.out1(R7134), .clock(clock), .in1(R7133));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7325 (.out1(R7326), .clock(clock), .in1(R7325));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7512 (.out1(R7513), .clock(clock), .in1(R7512));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7746 (.out1(R7747), .clock(clock), .in1(R7746));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7925 (.out1(R7926), .clock(clock), .in1(R7925));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8099 (.out1(R8100), .clock(clock), .in1(R8099));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8320 (.out1(R8321), .clock(clock), .in1(R8320));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8486 (.out1(R8487), .clock(clock), .in1(R8486));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8647 (.out1(R8648), .clock(clock), .in1(ifout611));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8815 (.out1(R8816), .clock(clock), .in1(_658));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8816 (.out1(R8817), .clock(clock), .in1(_651));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8817 (.out1(R8818), .clock(clock), .in1(_640));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8818 (.out1(R8819), .clock(clock), .in1(_620));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op654 (.out1(_632), .in1(R8321));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op634 (.out1(_612), .in1(R8321));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op623 (.out1(_601), .in1(R8321));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op616 (.out1(_594), .in1(R8321));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op683 (.out1(_661), .in1(2 'd 2), .in2(R8487));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op655 (.out1(_633), .in1(_632), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op635 (.out1(_613), .in1(_612), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op624 (.out1(_602), .in1(_601), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op617 (.out1(_595), .in1(_594), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op681 (.out1(_659), .in1(vec52_3587_D), .in2(R8816));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op674 (.out1(_652), .in1(vec52_3587_D), .in2(R8817));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op663 (.out1(_641), .in1(vec52_3587_D), .in2(R8818));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op643 (.out1(_621), .in1(vec52_3587_D), .in2(R8819));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3774 (.out1(R3775), .clock(clock), .in1(R3774));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4030 (.out1(R4031), .clock(clock), .in1(R4030));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4285 (.out1(R4286), .clock(clock), .in1(R4285));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4530 (.out1(R4531), .clock(clock), .in1(R4530));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4770 (.out1(R4771), .clock(clock), .in1(R4770));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5057 (.out1(R5058), .clock(clock), .in1(R5057));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5289 (.out1(R5290), .clock(clock), .in1(R5289));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5516 (.out1(R5517), .clock(clock), .in1(R5516));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5790 (.out1(R5791), .clock(clock), .in1(R5790));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6008 (.out1(R6009), .clock(clock), .in1(R6008));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6221 (.out1(R6222), .clock(clock), .in1(R6221));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6482 (.out1(R6483), .clock(clock), .in1(R6482));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6687 (.out1(R6688), .clock(clock), .in1(R6687));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6887 (.out1(R6888), .clock(clock), .in1(R6887));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7134 (.out1(R7135), .clock(clock), .in1(R7134));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7326 (.out1(R7327), .clock(clock), .in1(R7326));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7513 (.out1(R7514), .clock(clock), .in1(R7513));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7747 (.out1(R7748), .clock(clock), .in1(R7747));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7926 (.out1(R7927), .clock(clock), .in1(R7926));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8100 (.out1(R8101), .clock(clock), .in1(R8100));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8321 (.out1(R8322), .clock(clock), .in1(R8321));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8487 (.out1(R8488), .clock(clock), .in1(R8487));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8648 (.out1(R8649), .clock(clock), .in1(R8648));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8819 (.out1(R8820), .clock(clock), .in1(_661));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8820 (.out1(R8821), .clock(clock), .in1(_633));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8821 (.out1(R8822), .clock(clock), .in1(_613));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8822 (.out1(R8823), .clock(clock), .in1(_602));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8823 (.out1(R8824), .clock(clock), .in1(_595));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8824 (.out1(R8825), .clock(clock), .in1(_659));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8825 (.out1(R8826), .clock(clock), .in1(_652));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8826 (.out1(R8827), .clock(clock), .in1(_641));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8827 (.out1(R8828), .clock(clock), .in1(_621));
  SRAM op682 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_660),.ADR(R8825));
  SRAM op675 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_653),.ADR(R8826));
  SRAM op664 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_642),.ADR(R8827));
  SRAM op644 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_622),.ADR(R8828));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op676 (.out1(_654), .in1(2 'd 2), .in2(R8488));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op665 (.out1(_643), .in1(2 'd 2), .in2(R8488));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op658 (.out1(_636), .in1(2 'd 2), .in2(R8488));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op645 (.out1(_623), .in1(2 'd 2), .in2(R8488));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op638 (.out1(_616), .in1(2 'd 2), .in2(R8488));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op627 (.out1(_605), .in1(2 'd 2), .in2(R8488));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op656 (.out1(_634), .in1(vec52_3587_D), .in2(R8821));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op636 (.out1(_614), .in1(vec52_3587_D), .in2(R8822));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op625 (.out1(_603), .in1(vec52_3587_D), .in2(R8823));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op618 (.out1(_596), .in1(vec52_3587_D), .in2(R8824));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op684 (.out1(_662), .in1(R8820), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3775 (.out1(R3776), .clock(clock), .in1(R3775));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4031 (.out1(R4032), .clock(clock), .in1(R4031));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4286 (.out1(R4287), .clock(clock), .in1(R4286));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4531 (.out1(R4532), .clock(clock), .in1(R4531));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4771 (.out1(R4772), .clock(clock), .in1(R4771));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5058 (.out1(R5059), .clock(clock), .in1(R5058));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5290 (.out1(R5291), .clock(clock), .in1(R5290));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5517 (.out1(R5518), .clock(clock), .in1(R5517));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5791 (.out1(R5792), .clock(clock), .in1(R5791));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6009 (.out1(R6010), .clock(clock), .in1(R6009));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6222 (.out1(R6223), .clock(clock), .in1(R6222));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6483 (.out1(R6484), .clock(clock), .in1(R6483));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6688 (.out1(R6689), .clock(clock), .in1(R6688));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6888 (.out1(R6889), .clock(clock), .in1(R6888));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7135 (.out1(R7136), .clock(clock), .in1(R7135));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7327 (.out1(R7328), .clock(clock), .in1(R7327));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7514 (.out1(R7515), .clock(clock), .in1(R7514));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7748 (.out1(R7749), .clock(clock), .in1(R7748));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7927 (.out1(R7928), .clock(clock), .in1(R7927));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8101 (.out1(R8102), .clock(clock), .in1(R8101));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8322 (.out1(R8323), .clock(clock), .in1(R8322));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8488 (.out1(R8489), .clock(clock), .in1(R8488));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8649 (.out1(R8650), .clock(clock), .in1(R8649));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8828 (.out1(R8829), .clock(clock), .in1(_660));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8829 (.out1(R8830), .clock(clock), .in1(_653));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8830 (.out1(R8831), .clock(clock), .in1(_642));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8831 (.out1(R8832), .clock(clock), .in1(_622));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8832 (.out1(R8833), .clock(clock), .in1(_654));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8833 (.out1(R8834), .clock(clock), .in1(_643));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8834 (.out1(R8835), .clock(clock), .in1(_636));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8835 (.out1(R8836), .clock(clock), .in1(_623));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8836 (.out1(R8837), .clock(clock), .in1(_616));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8837 (.out1(R8838), .clock(clock), .in1(_605));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8838 (.out1(R8839), .clock(clock), .in1(_634));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8839 (.out1(R8840), .clock(clock), .in1(_614));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8840 (.out1(R8841), .clock(clock), .in1(_603));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8841 (.out1(R8842), .clock(clock), .in1(_596));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8842 (.out1(R8843), .clock(clock), .in1(_662));
  SRAM op657 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_635),.ADR(R8839));
  SRAM op637 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_615),.ADR(R8840));
  SRAM op626 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_604),.ADR(R8841));
  SRAM op619 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_597),.ADR(R8842));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op685 (.out1(_663), .in1(R8829), .in2(R8843));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op686 (.out1(_664), .in1(_663), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op677 (.out1(_655), .in1(R8833), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op666 (.out1(_644), .in1(R8834), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op646 (.out1(_624), .in1(R8836), .in2(64 'd 18446744073709551615));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op620 (.out1(_598), .in1(2 'd 2), .in2(R8489));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op687 (.out1(_665), .in1(_664), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op678 (.out1(_656), .in1(R8830), .in2(_655));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op667 (.out1(_645), .in1(R8831), .in2(_644));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op647 (.out1(_625), .in1(R8832), .in2(_624));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op688 (.out1(_666), .in1(_656), .in2(_665));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op668 (.out1(_646), .in1(_645), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op659 (.out1(_637), .in1(R8835), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op648 (.out1(_626), .in1(_625), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op639 (.out1(_617), .in1(R8837), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op628 (.out1(_606), .in1(R8838), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3776 (.out1(R3777), .clock(clock), .in1(R3776));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4032 (.out1(R4033), .clock(clock), .in1(R4032));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4287 (.out1(R4288), .clock(clock), .in1(R4287));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4532 (.out1(R4533), .clock(clock), .in1(R4532));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4772 (.out1(R4773), .clock(clock), .in1(R4772));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5059 (.out1(R5060), .clock(clock), .in1(R5059));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5291 (.out1(R5292), .clock(clock), .in1(R5291));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5518 (.out1(R5519), .clock(clock), .in1(R5518));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5792 (.out1(R5793), .clock(clock), .in1(R5792));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6010 (.out1(R6011), .clock(clock), .in1(R6010));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6223 (.out1(R6224), .clock(clock), .in1(R6223));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6484 (.out1(R6485), .clock(clock), .in1(R6484));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6689 (.out1(R6690), .clock(clock), .in1(R6689));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6889 (.out1(R6890), .clock(clock), .in1(R6889));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7136 (.out1(R7137), .clock(clock), .in1(R7136));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7328 (.out1(R7329), .clock(clock), .in1(R7328));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7515 (.out1(R7516), .clock(clock), .in1(R7515));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7749 (.out1(R7750), .clock(clock), .in1(R7749));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7928 (.out1(R7929), .clock(clock), .in1(R7928));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8102 (.out1(R8103), .clock(clock), .in1(R8102));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8323 (.out1(R8324), .clock(clock), .in1(R8323));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8489 (.out1(R8490), .clock(clock), .in1(R8489));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8650 (.out1(R8651), .clock(clock), .in1(R8650));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8843 (.out1(R8844), .clock(clock), .in1(_635));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8844 (.out1(R8845), .clock(clock), .in1(_615));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8845 (.out1(R8846), .clock(clock), .in1(_604));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8846 (.out1(R8847), .clock(clock), .in1(_597));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8847 (.out1(R8848), .clock(clock), .in1(_598));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8848 (.out1(R8849), .clock(clock), .in1(_666));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8849 (.out1(R8850), .clock(clock), .in1(_646));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8850 (.out1(R8851), .clock(clock), .in1(_637));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8851 (.out1(R8852), .clock(clock), .in1(_626));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8852 (.out1(R8853), .clock(clock), .in1(_617));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8853 (.out1(R8854), .clock(clock), .in1(_606));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op669 (.out1(_647), .in1(R8850), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op660 (.out1(_638), .in1(R8844), .in2(R8851));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op629 (.out1(_607), .in1(R8846), .in2(R8854));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op689 (.out1(_667), .in1(R8849), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op670 (.out1(_648), .in1(_638), .in2(_647));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op649 (.out1(_627), .in1(R8852), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op640 (.out1(_618), .in1(R8845), .in2(R8853));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op630 (.out1(_608), .in1(_607), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op621 (.out1(_599), .in1(R8848), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op650 (.out1(_628), .in1(_618), .in2(_627));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op690 (.out1(_668), .in1(_667), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op671 (.out1(_649), .in1(_648), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op631 (.out1(_609), .in1(_608), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op622 (.out1(_600), .in1(R8847), .in2(_599));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op691 (.out1(_669), .in1(_649), .in2(_668));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op651 (.out1(_629), .in1(_628), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op632 (.out1(_610), .in1(_600), .in2(_609));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3777 (.out1(R3778), .clock(clock), .in1(R3777));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4033 (.out1(R4034), .clock(clock), .in1(R4033));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4288 (.out1(R4289), .clock(clock), .in1(R4288));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4533 (.out1(R4534), .clock(clock), .in1(R4533));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4773 (.out1(R4774), .clock(clock), .in1(R4773));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5060 (.out1(R5061), .clock(clock), .in1(R5060));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5292 (.out1(R5293), .clock(clock), .in1(R5292));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5519 (.out1(R5520), .clock(clock), .in1(R5519));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5793 (.out1(R5794), .clock(clock), .in1(R5793));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6011 (.out1(R6012), .clock(clock), .in1(R6011));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6224 (.out1(R6225), .clock(clock), .in1(R6224));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6485 (.out1(R6486), .clock(clock), .in1(R6485));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6690 (.out1(R6691), .clock(clock), .in1(R6690));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6890 (.out1(R6891), .clock(clock), .in1(R6890));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7137 (.out1(R7138), .clock(clock), .in1(R7137));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7329 (.out1(R7330), .clock(clock), .in1(R7329));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7516 (.out1(R7517), .clock(clock), .in1(R7516));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7750 (.out1(R7751), .clock(clock), .in1(R7750));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7929 (.out1(R7930), .clock(clock), .in1(R7929));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8103 (.out1(R8104), .clock(clock), .in1(R8103));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8324 (.out1(R8325), .clock(clock), .in1(R8324));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8490 (.out1(R8491), .clock(clock), .in1(R8490));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8651 (.out1(R8652), .clock(clock), .in1(R8651));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8854 (.out1(R8855), .clock(clock), .in1(_669));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8855 (.out1(R8856), .clock(clock), .in1(_629));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8856 (.out1(R8857), .clock(clock), .in1(_610));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op612 (.out1(_590), .in1(R8325));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op652 (.out1(_630), .in1(R8856), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op633 (.out1(_611), .in1(R8857), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op692 (.out1(_670), .in1(R8855), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op653 (.out1(_631), .in1(_611), .in2(_630));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op613 (.out1(_591), .in1(_590), .in2(2 'd 2));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op693 (.out1(_671), .in1(_631), .in2(_670));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op694 (.out1(_672), .in1(_671), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3778 (.out1(R3779), .clock(clock), .in1(R3778));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4034 (.out1(R4035), .clock(clock), .in1(R4034));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4289 (.out1(R4290), .clock(clock), .in1(R4289));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4534 (.out1(R4535), .clock(clock), .in1(R4534));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4774 (.out1(R4775), .clock(clock), .in1(R4774));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5061 (.out1(R5062), .clock(clock), .in1(R5061));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5293 (.out1(R5294), .clock(clock), .in1(R5293));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5520 (.out1(R5521), .clock(clock), .in1(R5520));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5794 (.out1(R5795), .clock(clock), .in1(R5794));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6012 (.out1(R6013), .clock(clock), .in1(R6012));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6225 (.out1(R6226), .clock(clock), .in1(R6225));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6486 (.out1(R6487), .clock(clock), .in1(R6486));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6691 (.out1(R6692), .clock(clock), .in1(R6691));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6891 (.out1(R6892), .clock(clock), .in1(R6891));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7138 (.out1(R7139), .clock(clock), .in1(R7138));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7330 (.out1(R7331), .clock(clock), .in1(R7330));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7517 (.out1(R7518), .clock(clock), .in1(R7517));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7751 (.out1(R7752), .clock(clock), .in1(R7751));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7930 (.out1(R7931), .clock(clock), .in1(R7930));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8104 (.out1(R8105), .clock(clock), .in1(R8104));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8325 (.out1(R8326), .clock(clock), .in1(R8325));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8491 (.out1(R8492), .clock(clock), .in1(R8491));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8652 (.out1(R8653), .clock(clock), .in1(R8652));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8857 (.out1(R8858), .clock(clock), .in1(_591));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8858 (.out1(R8859), .clock(clock), .in1(_672));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op695 (.out1(_673), .in1(R8859), .in2(57 'd 72340172838076673));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op614 (.out1(_592), .in1(base0_52_3592_D), .in2(R8858));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3779 (.out1(R3780), .clock(clock), .in1(R3779));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4035 (.out1(R4036), .clock(clock), .in1(R4035));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4290 (.out1(R4291), .clock(clock), .in1(R4290));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4535 (.out1(R4536), .clock(clock), .in1(R4535));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4775 (.out1(R4776), .clock(clock), .in1(R4775));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5062 (.out1(R5063), .clock(clock), .in1(R5062));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5294 (.out1(R5295), .clock(clock), .in1(R5294));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5521 (.out1(R5522), .clock(clock), .in1(R5521));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5795 (.out1(R5796), .clock(clock), .in1(R5795));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6013 (.out1(R6014), .clock(clock), .in1(R6013));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6226 (.out1(R6227), .clock(clock), .in1(R6226));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6487 (.out1(R6488), .clock(clock), .in1(R6487));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6692 (.out1(R6693), .clock(clock), .in1(R6692));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6892 (.out1(R6893), .clock(clock), .in1(R6892));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7139 (.out1(R7140), .clock(clock), .in1(R7139));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7331 (.out1(R7332), .clock(clock), .in1(R7331));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7518 (.out1(R7519), .clock(clock), .in1(R7518));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7752 (.out1(R7753), .clock(clock), .in1(R7752));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7931 (.out1(R7932), .clock(clock), .in1(R7931));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8105 (.out1(R8106), .clock(clock), .in1(R8105));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8326 (.out1(R8327), .clock(clock), .in1(R8326));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8492 (.out1(R8493), .clock(clock), .in1(R8492));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8653 (.out1(R8654), .clock(clock), .in1(R8653));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8859 (.out1(R8860), .clock(clock), .in1(_673));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8860 (.out1(R8861), .clock(clock), .in1(_592));
  SRAM op615 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_593),.ADR(R8861));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op696 (.out1(_674), .in1(R8860), .in2(6 'd 56));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3780 (.out1(R3781), .clock(clock), .in1(R3780));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4036 (.out1(R4037), .clock(clock), .in1(R4036));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4291 (.out1(R4292), .clock(clock), .in1(R4291));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4536 (.out1(R4537), .clock(clock), .in1(R4536));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4776 (.out1(R4777), .clock(clock), .in1(R4776));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5063 (.out1(R5064), .clock(clock), .in1(R5063));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5295 (.out1(R5296), .clock(clock), .in1(R5295));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5522 (.out1(R5523), .clock(clock), .in1(R5522));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5796 (.out1(R5797), .clock(clock), .in1(R5796));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6014 (.out1(R6015), .clock(clock), .in1(R6014));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6227 (.out1(R6228), .clock(clock), .in1(R6227));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6488 (.out1(R6489), .clock(clock), .in1(R6488));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6693 (.out1(R6694), .clock(clock), .in1(R6693));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6893 (.out1(R6894), .clock(clock), .in1(R6893));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7140 (.out1(R7141), .clock(clock), .in1(R7140));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7332 (.out1(R7333), .clock(clock), .in1(R7332));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7519 (.out1(R7520), .clock(clock), .in1(R7519));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7753 (.out1(R7754), .clock(clock), .in1(R7753));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7932 (.out1(R7933), .clock(clock), .in1(R7932));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8106 (.out1(R8107), .clock(clock), .in1(R8106));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8327 (.out1(R8328), .clock(clock), .in1(R8327));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8493 (.out1(R8494), .clock(clock), .in1(R8493));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8654 (.out1(R8655), .clock(clock), .in1(R8654));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8861 (.out1(R8862), .clock(clock), .in1(_593));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op8862 (.out1(R8863), .clock(clock), .in1(_674));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op697 (.out1(_675), .in1(R8863));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op698 (.out1(_676), .in1(R8862), .in2(_675));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op699 (.out1(idx_3593), .in1(_676), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3781 (.out1(R3782), .clock(clock), .in1(R3781));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4037 (.out1(R4038), .clock(clock), .in1(R4037));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4292 (.out1(R4293), .clock(clock), .in1(R4292));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4537 (.out1(R4538), .clock(clock), .in1(R4537));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4777 (.out1(R4778), .clock(clock), .in1(R4777));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5064 (.out1(R5065), .clock(clock), .in1(R5064));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5296 (.out1(R5297), .clock(clock), .in1(R5296));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5523 (.out1(R5524), .clock(clock), .in1(R5523));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5797 (.out1(R5798), .clock(clock), .in1(R5797));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6015 (.out1(R6016), .clock(clock), .in1(R6015));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6228 (.out1(R6229), .clock(clock), .in1(R6228));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6489 (.out1(R6490), .clock(clock), .in1(R6489));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6694 (.out1(R6695), .clock(clock), .in1(R6694));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6894 (.out1(R6895), .clock(clock), .in1(R6894));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7141 (.out1(R7142), .clock(clock), .in1(R7141));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7333 (.out1(R7334), .clock(clock), .in1(R7333));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7520 (.out1(R7521), .clock(clock), .in1(R7520));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7754 (.out1(R7755), .clock(clock), .in1(R7754));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7933 (.out1(R7934), .clock(clock), .in1(R7933));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8107 (.out1(R8108), .clock(clock), .in1(R8107));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8328 (.out1(R8329), .clock(clock), .in1(R8328));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8494 (.out1(R8495), .clock(clock), .in1(R8494));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8655 (.out1(R8656), .clock(clock), .in1(R8655));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8863 (.out1(R8864), .clock(clock), .in1(idx_3593));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op702 (.out1(_678), .in1(R8864));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op703 (.out1(_679), .in1(_678), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3782 (.out1(R3783), .clock(clock), .in1(R3782));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4038 (.out1(R4039), .clock(clock), .in1(R4038));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4293 (.out1(R4294), .clock(clock), .in1(R4293));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4538 (.out1(R4539), .clock(clock), .in1(R4538));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4778 (.out1(R4779), .clock(clock), .in1(R4778));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5065 (.out1(R5066), .clock(clock), .in1(R5065));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5297 (.out1(R5298), .clock(clock), .in1(R5297));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5524 (.out1(R5525), .clock(clock), .in1(R5524));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5798 (.out1(R5799), .clock(clock), .in1(R5798));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6016 (.out1(R6017), .clock(clock), .in1(R6016));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6229 (.out1(R6230), .clock(clock), .in1(R6229));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6490 (.out1(R6491), .clock(clock), .in1(R6490));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6695 (.out1(R6696), .clock(clock), .in1(R6695));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6895 (.out1(R6896), .clock(clock), .in1(R6895));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7142 (.out1(R7143), .clock(clock), .in1(R7142));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7334 (.out1(R7335), .clock(clock), .in1(R7334));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7521 (.out1(R7522), .clock(clock), .in1(R7521));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7755 (.out1(R7756), .clock(clock), .in1(R7755));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7934 (.out1(R7935), .clock(clock), .in1(R7934));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8108 (.out1(R8109), .clock(clock), .in1(R8108));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8329 (.out1(R8330), .clock(clock), .in1(R8329));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8495 (.out1(R8496), .clock(clock), .in1(R8495));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8656 (.out1(R8657), .clock(clock), .in1(R8656));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8864 (.out1(R8865), .clock(clock), .in1(R8864));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9017 (.out1(R9018), .clock(clock), .in1(_679));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op704 (.out1(_680), .in1(vec58_3595_D), .in2(R9018));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3783 (.out1(R3784), .clock(clock), .in1(R3783));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4039 (.out1(R4040), .clock(clock), .in1(R4039));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4294 (.out1(R4295), .clock(clock), .in1(R4294));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4539 (.out1(R4540), .clock(clock), .in1(R4539));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4779 (.out1(R4780), .clock(clock), .in1(R4779));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5066 (.out1(R5067), .clock(clock), .in1(R5066));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5298 (.out1(R5299), .clock(clock), .in1(R5298));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5525 (.out1(R5526), .clock(clock), .in1(R5525));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5799 (.out1(R5800), .clock(clock), .in1(R5799));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6017 (.out1(R6018), .clock(clock), .in1(R6017));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6230 (.out1(R6231), .clock(clock), .in1(R6230));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6491 (.out1(R6492), .clock(clock), .in1(R6491));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6696 (.out1(R6697), .clock(clock), .in1(R6696));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6896 (.out1(R6897), .clock(clock), .in1(R6896));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7143 (.out1(R7144), .clock(clock), .in1(R7143));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7335 (.out1(R7336), .clock(clock), .in1(R7335));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7522 (.out1(R7523), .clock(clock), .in1(R7522));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7756 (.out1(R7757), .clock(clock), .in1(R7756));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7935 (.out1(R7936), .clock(clock), .in1(R7935));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8109 (.out1(R8110), .clock(clock), .in1(R8109));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8330 (.out1(R8331), .clock(clock), .in1(R8330));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8496 (.out1(R8497), .clock(clock), .in1(R8496));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8657 (.out1(R8658), .clock(clock), .in1(R8657));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8865 (.out1(R8866), .clock(clock), .in1(R8865));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9018 (.out1(R9019), .clock(clock), .in1(_680));
  SRAM op705 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_681),.ADR(R9019));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3784 (.out1(R3785), .clock(clock), .in1(R3784));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4040 (.out1(R4041), .clock(clock), .in1(R4040));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4295 (.out1(R4296), .clock(clock), .in1(R4295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4540 (.out1(R4541), .clock(clock), .in1(R4540));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4780 (.out1(R4781), .clock(clock), .in1(R4780));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5067 (.out1(R5068), .clock(clock), .in1(R5067));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5299 (.out1(R5300), .clock(clock), .in1(R5299));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5526 (.out1(R5527), .clock(clock), .in1(R5526));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5800 (.out1(R5801), .clock(clock), .in1(R5800));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6018 (.out1(R6019), .clock(clock), .in1(R6018));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6231 (.out1(R6232), .clock(clock), .in1(R6231));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6492 (.out1(R6493), .clock(clock), .in1(R6492));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6697 (.out1(R6698), .clock(clock), .in1(R6697));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6897 (.out1(R6898), .clock(clock), .in1(R6897));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7144 (.out1(R7145), .clock(clock), .in1(R7144));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7336 (.out1(R7337), .clock(clock), .in1(R7336));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7523 (.out1(R7524), .clock(clock), .in1(R7523));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7757 (.out1(R7758), .clock(clock), .in1(R7757));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7936 (.out1(R7937), .clock(clock), .in1(R7936));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8110 (.out1(R8111), .clock(clock), .in1(R8110));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8331 (.out1(R8332), .clock(clock), .in1(R8331));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8497 (.out1(R8498), .clock(clock), .in1(R8497));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8658 (.out1(R8659), .clock(clock), .in1(R8658));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8866 (.out1(R8867), .clock(clock), .in1(R8866));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9019 (.out1(R9020), .clock(clock), .in1(_681));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op700 (.out1(_677), .in1(ip1_3530_D));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op701 (.out1(off_3594), .in1(_677), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op706 (.out1(_682), .in1(R9020), .in2(off_3594));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3785 (.out1(R3786), .clock(clock), .in1(R3785));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4041 (.out1(R4042), .clock(clock), .in1(R4041));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4296 (.out1(R4297), .clock(clock), .in1(R4296));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4541 (.out1(R4542), .clock(clock), .in1(R4541));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4781 (.out1(R4782), .clock(clock), .in1(R4781));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5068 (.out1(R5069), .clock(clock), .in1(R5068));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5300 (.out1(R5301), .clock(clock), .in1(R5300));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5527 (.out1(R5528), .clock(clock), .in1(R5527));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5801 (.out1(R5802), .clock(clock), .in1(R5801));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6019 (.out1(R6020), .clock(clock), .in1(R6019));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6232 (.out1(R6233), .clock(clock), .in1(R6232));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6493 (.out1(R6494), .clock(clock), .in1(R6493));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6698 (.out1(R6699), .clock(clock), .in1(R6698));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6898 (.out1(R6899), .clock(clock), .in1(R6898));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7145 (.out1(R7146), .clock(clock), .in1(R7145));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7337 (.out1(R7338), .clock(clock), .in1(R7337));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7524 (.out1(R7525), .clock(clock), .in1(R7524));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7758 (.out1(R7759), .clock(clock), .in1(R7758));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7937 (.out1(R7938), .clock(clock), .in1(R7937));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8111 (.out1(R8112), .clock(clock), .in1(R8111));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8332 (.out1(R8333), .clock(clock), .in1(R8332));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8498 (.out1(R8499), .clock(clock), .in1(R8498));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8659 (.out1(R8660), .clock(clock), .in1(R8659));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8867 (.out1(R8868), .clock(clock), .in1(R8867));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9020 (.out1(R9021), .clock(clock), .in1(off_3594));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9168 (.out1(R9169), .clock(clock), .in1(_682));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op707 (.out1(_683), .in1(R9169), .in2(1 'd 1));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op708 (.out1(ifout708), .in1(_683), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op776 (.out1(_751), .in1(R8868));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op769 (.out1(_744), .in1(R8868));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op758 (.out1(_733), .in1(R8868));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op738 (.out1(_713), .in1(R8868));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op777 (.out1(_752), .in1(_751), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op770 (.out1(_745), .in1(_744), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op759 (.out1(_734), .in1(_733), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op739 (.out1(_714), .in1(_713), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3786 (.out1(R3787), .clock(clock), .in1(R3786));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4042 (.out1(R4043), .clock(clock), .in1(R4042));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4297 (.out1(R4298), .clock(clock), .in1(R4297));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4542 (.out1(R4543), .clock(clock), .in1(R4542));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4782 (.out1(R4783), .clock(clock), .in1(R4782));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5069 (.out1(R5070), .clock(clock), .in1(R5069));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5301 (.out1(R5302), .clock(clock), .in1(R5301));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5528 (.out1(R5529), .clock(clock), .in1(R5528));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5802 (.out1(R5803), .clock(clock), .in1(R5802));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6020 (.out1(R6021), .clock(clock), .in1(R6020));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6233 (.out1(R6234), .clock(clock), .in1(R6233));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6494 (.out1(R6495), .clock(clock), .in1(R6494));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6699 (.out1(R6700), .clock(clock), .in1(R6699));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6899 (.out1(R6900), .clock(clock), .in1(R6899));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7146 (.out1(R7147), .clock(clock), .in1(R7146));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7338 (.out1(R7339), .clock(clock), .in1(R7338));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7525 (.out1(R7526), .clock(clock), .in1(R7525));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7759 (.out1(R7760), .clock(clock), .in1(R7759));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7938 (.out1(R7939), .clock(clock), .in1(R7938));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8112 (.out1(R8113), .clock(clock), .in1(R8112));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8333 (.out1(R8334), .clock(clock), .in1(R8333));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8499 (.out1(R8500), .clock(clock), .in1(R8499));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8660 (.out1(R8661), .clock(clock), .in1(R8660));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8868 (.out1(R8869), .clock(clock), .in1(R8868));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9021 (.out1(R9022), .clock(clock), .in1(R9021));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9169 (.out1(R9170), .clock(clock), .in1(ifout708));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9324 (.out1(R9325), .clock(clock), .in1(_752));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9325 (.out1(R9326), .clock(clock), .in1(_745));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9326 (.out1(R9327), .clock(clock), .in1(_734));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9327 (.out1(R9328), .clock(clock), .in1(_714));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op751 (.out1(_726), .in1(R8869));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op731 (.out1(_706), .in1(R8869));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op720 (.out1(_695), .in1(R8869));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op713 (.out1(_688), .in1(R8869));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op780 (.out1(_755), .in1(2 'd 2), .in2(R9022));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op752 (.out1(_727), .in1(_726), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op732 (.out1(_707), .in1(_706), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op721 (.out1(_696), .in1(_695), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op714 (.out1(_689), .in1(_688), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op778 (.out1(_753), .in1(vec58_3595_D), .in2(R9325));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op771 (.out1(_746), .in1(vec58_3595_D), .in2(R9326));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op760 (.out1(_735), .in1(vec58_3595_D), .in2(R9327));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op740 (.out1(_715), .in1(vec58_3595_D), .in2(R9328));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3787 (.out1(R3788), .clock(clock), .in1(R3787));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4043 (.out1(R4044), .clock(clock), .in1(R4043));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4298 (.out1(R4299), .clock(clock), .in1(R4298));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4543 (.out1(R4544), .clock(clock), .in1(R4543));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4783 (.out1(R4784), .clock(clock), .in1(R4783));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5070 (.out1(R5071), .clock(clock), .in1(R5070));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5302 (.out1(R5303), .clock(clock), .in1(R5302));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5529 (.out1(R5530), .clock(clock), .in1(R5529));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5803 (.out1(R5804), .clock(clock), .in1(R5803));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6021 (.out1(R6022), .clock(clock), .in1(R6021));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6234 (.out1(R6235), .clock(clock), .in1(R6234));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6495 (.out1(R6496), .clock(clock), .in1(R6495));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6700 (.out1(R6701), .clock(clock), .in1(R6700));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6900 (.out1(R6901), .clock(clock), .in1(R6900));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7147 (.out1(R7148), .clock(clock), .in1(R7147));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7339 (.out1(R7340), .clock(clock), .in1(R7339));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7526 (.out1(R7527), .clock(clock), .in1(R7526));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7760 (.out1(R7761), .clock(clock), .in1(R7760));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7939 (.out1(R7940), .clock(clock), .in1(R7939));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8113 (.out1(R8114), .clock(clock), .in1(R8113));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8334 (.out1(R8335), .clock(clock), .in1(R8334));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8500 (.out1(R8501), .clock(clock), .in1(R8500));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8661 (.out1(R8662), .clock(clock), .in1(R8661));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8869 (.out1(R8870), .clock(clock), .in1(R8869));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9022 (.out1(R9023), .clock(clock), .in1(R9022));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9170 (.out1(R9171), .clock(clock), .in1(R9170));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9328 (.out1(R9329), .clock(clock), .in1(_755));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9329 (.out1(R9330), .clock(clock), .in1(_727));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9330 (.out1(R9331), .clock(clock), .in1(_707));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9331 (.out1(R9332), .clock(clock), .in1(_696));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9332 (.out1(R9333), .clock(clock), .in1(_689));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9333 (.out1(R9334), .clock(clock), .in1(_753));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9334 (.out1(R9335), .clock(clock), .in1(_746));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9335 (.out1(R9336), .clock(clock), .in1(_735));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9336 (.out1(R9337), .clock(clock), .in1(_715));
  SRAM op779 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_754),.ADR(R9334));
  SRAM op772 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_747),.ADR(R9335));
  SRAM op761 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_736),.ADR(R9336));
  SRAM op741 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_716),.ADR(R9337));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op773 (.out1(_748), .in1(2 'd 2), .in2(R9023));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op762 (.out1(_737), .in1(2 'd 2), .in2(R9023));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op755 (.out1(_730), .in1(2 'd 2), .in2(R9023));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op742 (.out1(_717), .in1(2 'd 2), .in2(R9023));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op735 (.out1(_710), .in1(2 'd 2), .in2(R9023));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op724 (.out1(_699), .in1(2 'd 2), .in2(R9023));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op753 (.out1(_728), .in1(vec58_3595_D), .in2(R9330));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op733 (.out1(_708), .in1(vec58_3595_D), .in2(R9331));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op722 (.out1(_697), .in1(vec58_3595_D), .in2(R9332));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op715 (.out1(_690), .in1(vec58_3595_D), .in2(R9333));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op781 (.out1(_756), .in1(R9329), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3788 (.out1(R3789), .clock(clock), .in1(R3788));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4044 (.out1(R4045), .clock(clock), .in1(R4044));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4299 (.out1(R4300), .clock(clock), .in1(R4299));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4544 (.out1(R4545), .clock(clock), .in1(R4544));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4784 (.out1(R4785), .clock(clock), .in1(R4784));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5071 (.out1(R5072), .clock(clock), .in1(R5071));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5303 (.out1(R5304), .clock(clock), .in1(R5303));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5530 (.out1(R5531), .clock(clock), .in1(R5530));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5804 (.out1(R5805), .clock(clock), .in1(R5804));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6022 (.out1(R6023), .clock(clock), .in1(R6022));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6235 (.out1(R6236), .clock(clock), .in1(R6235));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6496 (.out1(R6497), .clock(clock), .in1(R6496));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6701 (.out1(R6702), .clock(clock), .in1(R6701));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6901 (.out1(R6902), .clock(clock), .in1(R6901));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7148 (.out1(R7149), .clock(clock), .in1(R7148));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7340 (.out1(R7341), .clock(clock), .in1(R7340));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7527 (.out1(R7528), .clock(clock), .in1(R7527));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7761 (.out1(R7762), .clock(clock), .in1(R7761));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7940 (.out1(R7941), .clock(clock), .in1(R7940));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8114 (.out1(R8115), .clock(clock), .in1(R8114));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8335 (.out1(R8336), .clock(clock), .in1(R8335));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8501 (.out1(R8502), .clock(clock), .in1(R8501));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8662 (.out1(R8663), .clock(clock), .in1(R8662));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8870 (.out1(R8871), .clock(clock), .in1(R8870));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9023 (.out1(R9024), .clock(clock), .in1(R9023));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9171 (.out1(R9172), .clock(clock), .in1(R9171));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9337 (.out1(R9338), .clock(clock), .in1(_754));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9338 (.out1(R9339), .clock(clock), .in1(_747));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9339 (.out1(R9340), .clock(clock), .in1(_736));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9340 (.out1(R9341), .clock(clock), .in1(_716));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9341 (.out1(R9342), .clock(clock), .in1(_748));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9342 (.out1(R9343), .clock(clock), .in1(_737));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9343 (.out1(R9344), .clock(clock), .in1(_730));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9344 (.out1(R9345), .clock(clock), .in1(_717));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9345 (.out1(R9346), .clock(clock), .in1(_710));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9346 (.out1(R9347), .clock(clock), .in1(_699));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9347 (.out1(R9348), .clock(clock), .in1(_728));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9348 (.out1(R9349), .clock(clock), .in1(_708));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9349 (.out1(R9350), .clock(clock), .in1(_697));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9350 (.out1(R9351), .clock(clock), .in1(_690));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9351 (.out1(R9352), .clock(clock), .in1(_756));
  SRAM op754 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_729),.ADR(R9348));
  SRAM op734 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_709),.ADR(R9349));
  SRAM op723 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_698),.ADR(R9350));
  SRAM op716 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_691),.ADR(R9351));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op782 (.out1(_757), .in1(R9338), .in2(R9352));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op783 (.out1(_758), .in1(_757), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op774 (.out1(_749), .in1(R9342), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op763 (.out1(_738), .in1(R9343), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op743 (.out1(_718), .in1(R9345), .in2(64 'd 18446744073709551615));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op717 (.out1(_692), .in1(2 'd 2), .in2(R9024));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op784 (.out1(_759), .in1(_758), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op775 (.out1(_750), .in1(R9339), .in2(_749));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op764 (.out1(_739), .in1(R9340), .in2(_738));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op744 (.out1(_719), .in1(R9341), .in2(_718));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op785 (.out1(_760), .in1(_750), .in2(_759));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op765 (.out1(_740), .in1(_739), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op756 (.out1(_731), .in1(R9344), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op745 (.out1(_720), .in1(_719), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op736 (.out1(_711), .in1(R9346), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op725 (.out1(_700), .in1(R9347), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3789 (.out1(R3790), .clock(clock), .in1(R3789));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4045 (.out1(R4046), .clock(clock), .in1(R4045));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4300 (.out1(R4301), .clock(clock), .in1(R4300));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4545 (.out1(R4546), .clock(clock), .in1(R4545));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4785 (.out1(R4786), .clock(clock), .in1(R4785));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5072 (.out1(R5073), .clock(clock), .in1(R5072));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5304 (.out1(R5305), .clock(clock), .in1(R5304));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5531 (.out1(R5532), .clock(clock), .in1(R5531));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5805 (.out1(R5806), .clock(clock), .in1(R5805));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6023 (.out1(R6024), .clock(clock), .in1(R6023));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6236 (.out1(R6237), .clock(clock), .in1(R6236));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6497 (.out1(R6498), .clock(clock), .in1(R6497));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6702 (.out1(R6703), .clock(clock), .in1(R6702));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6902 (.out1(R6903), .clock(clock), .in1(R6902));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7149 (.out1(R7150), .clock(clock), .in1(R7149));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7341 (.out1(R7342), .clock(clock), .in1(R7341));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7528 (.out1(R7529), .clock(clock), .in1(R7528));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7762 (.out1(R7763), .clock(clock), .in1(R7762));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7941 (.out1(R7942), .clock(clock), .in1(R7941));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8115 (.out1(R8116), .clock(clock), .in1(R8115));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8336 (.out1(R8337), .clock(clock), .in1(R8336));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8502 (.out1(R8503), .clock(clock), .in1(R8502));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8663 (.out1(R8664), .clock(clock), .in1(R8663));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8871 (.out1(R8872), .clock(clock), .in1(R8871));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9024 (.out1(R9025), .clock(clock), .in1(R9024));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9172 (.out1(R9173), .clock(clock), .in1(R9172));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9352 (.out1(R9353), .clock(clock), .in1(_729));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9353 (.out1(R9354), .clock(clock), .in1(_709));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9354 (.out1(R9355), .clock(clock), .in1(_698));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9355 (.out1(R9356), .clock(clock), .in1(_691));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9356 (.out1(R9357), .clock(clock), .in1(_692));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9357 (.out1(R9358), .clock(clock), .in1(_760));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9358 (.out1(R9359), .clock(clock), .in1(_740));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9359 (.out1(R9360), .clock(clock), .in1(_731));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9360 (.out1(R9361), .clock(clock), .in1(_720));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9361 (.out1(R9362), .clock(clock), .in1(_711));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9362 (.out1(R9363), .clock(clock), .in1(_700));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op766 (.out1(_741), .in1(R9359), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op757 (.out1(_732), .in1(R9353), .in2(R9360));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op726 (.out1(_701), .in1(R9355), .in2(R9363));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op786 (.out1(_761), .in1(R9358), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op767 (.out1(_742), .in1(_732), .in2(_741));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op746 (.out1(_721), .in1(R9361), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op737 (.out1(_712), .in1(R9354), .in2(R9362));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op727 (.out1(_702), .in1(_701), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op718 (.out1(_693), .in1(R9357), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op747 (.out1(_722), .in1(_712), .in2(_721));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op787 (.out1(_762), .in1(_761), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op768 (.out1(_743), .in1(_742), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op728 (.out1(_703), .in1(_702), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op719 (.out1(_694), .in1(R9356), .in2(_693));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op788 (.out1(_763), .in1(_743), .in2(_762));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op748 (.out1(_723), .in1(_722), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op729 (.out1(_704), .in1(_694), .in2(_703));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3790 (.out1(R3791), .clock(clock), .in1(R3790));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4046 (.out1(R4047), .clock(clock), .in1(R4046));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4301 (.out1(R4302), .clock(clock), .in1(R4301));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4546 (.out1(R4547), .clock(clock), .in1(R4546));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4786 (.out1(R4787), .clock(clock), .in1(R4786));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5073 (.out1(R5074), .clock(clock), .in1(R5073));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5305 (.out1(R5306), .clock(clock), .in1(R5305));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5532 (.out1(R5533), .clock(clock), .in1(R5532));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5806 (.out1(R5807), .clock(clock), .in1(R5806));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6024 (.out1(R6025), .clock(clock), .in1(R6024));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6237 (.out1(R6238), .clock(clock), .in1(R6237));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6498 (.out1(R6499), .clock(clock), .in1(R6498));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6703 (.out1(R6704), .clock(clock), .in1(R6703));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6903 (.out1(R6904), .clock(clock), .in1(R6903));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7150 (.out1(R7151), .clock(clock), .in1(R7150));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7342 (.out1(R7343), .clock(clock), .in1(R7342));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7529 (.out1(R7530), .clock(clock), .in1(R7529));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7763 (.out1(R7764), .clock(clock), .in1(R7763));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7942 (.out1(R7943), .clock(clock), .in1(R7942));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8116 (.out1(R8117), .clock(clock), .in1(R8116));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8337 (.out1(R8338), .clock(clock), .in1(R8337));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8503 (.out1(R8504), .clock(clock), .in1(R8503));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8664 (.out1(R8665), .clock(clock), .in1(R8664));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8872 (.out1(R8873), .clock(clock), .in1(R8872));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9025 (.out1(R9026), .clock(clock), .in1(R9025));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9173 (.out1(R9174), .clock(clock), .in1(R9173));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9363 (.out1(R9364), .clock(clock), .in1(_763));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9364 (.out1(R9365), .clock(clock), .in1(_723));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9365 (.out1(R9366), .clock(clock), .in1(_704));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op709 (.out1(_684), .in1(R8873));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op749 (.out1(_724), .in1(R9365), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op730 (.out1(_705), .in1(R9366), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op789 (.out1(_764), .in1(R9364), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op750 (.out1(_725), .in1(_705), .in2(_724));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op710 (.out1(_685), .in1(_684), .in2(2 'd 2));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op790 (.out1(_765), .in1(_725), .in2(_764));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op791 (.out1(_766), .in1(_765), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3791 (.out1(R3792), .clock(clock), .in1(R3791));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4047 (.out1(R4048), .clock(clock), .in1(R4047));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4302 (.out1(R4303), .clock(clock), .in1(R4302));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4547 (.out1(R4548), .clock(clock), .in1(R4547));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4787 (.out1(R4788), .clock(clock), .in1(R4787));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5074 (.out1(R5075), .clock(clock), .in1(R5074));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5306 (.out1(R5307), .clock(clock), .in1(R5306));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5533 (.out1(R5534), .clock(clock), .in1(R5533));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5807 (.out1(R5808), .clock(clock), .in1(R5807));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6025 (.out1(R6026), .clock(clock), .in1(R6025));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6238 (.out1(R6239), .clock(clock), .in1(R6238));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6499 (.out1(R6500), .clock(clock), .in1(R6499));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6704 (.out1(R6705), .clock(clock), .in1(R6704));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6904 (.out1(R6905), .clock(clock), .in1(R6904));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7151 (.out1(R7152), .clock(clock), .in1(R7151));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7343 (.out1(R7344), .clock(clock), .in1(R7343));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7530 (.out1(R7531), .clock(clock), .in1(R7530));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7764 (.out1(R7765), .clock(clock), .in1(R7764));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7943 (.out1(R7944), .clock(clock), .in1(R7943));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8117 (.out1(R8118), .clock(clock), .in1(R8117));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8338 (.out1(R8339), .clock(clock), .in1(R8338));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8504 (.out1(R8505), .clock(clock), .in1(R8504));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8665 (.out1(R8666), .clock(clock), .in1(R8665));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8873 (.out1(R8874), .clock(clock), .in1(R8873));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9026 (.out1(R9027), .clock(clock), .in1(R9026));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9174 (.out1(R9175), .clock(clock), .in1(R9174));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9366 (.out1(R9367), .clock(clock), .in1(_685));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9367 (.out1(R9368), .clock(clock), .in1(_766));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op792 (.out1(_767), .in1(R9368), .in2(57 'd 72340172838076673));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op711 (.out1(_686), .in1(base0_58_3600_D), .in2(R9367));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3792 (.out1(R3793), .clock(clock), .in1(R3792));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4048 (.out1(R4049), .clock(clock), .in1(R4048));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4303 (.out1(R4304), .clock(clock), .in1(R4303));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4548 (.out1(R4549), .clock(clock), .in1(R4548));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4788 (.out1(R4789), .clock(clock), .in1(R4788));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5075 (.out1(R5076), .clock(clock), .in1(R5075));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5307 (.out1(R5308), .clock(clock), .in1(R5307));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5534 (.out1(R5535), .clock(clock), .in1(R5534));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5808 (.out1(R5809), .clock(clock), .in1(R5808));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6026 (.out1(R6027), .clock(clock), .in1(R6026));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6239 (.out1(R6240), .clock(clock), .in1(R6239));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6500 (.out1(R6501), .clock(clock), .in1(R6500));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6705 (.out1(R6706), .clock(clock), .in1(R6705));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6905 (.out1(R6906), .clock(clock), .in1(R6905));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7152 (.out1(R7153), .clock(clock), .in1(R7152));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7344 (.out1(R7345), .clock(clock), .in1(R7344));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7531 (.out1(R7532), .clock(clock), .in1(R7531));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7765 (.out1(R7766), .clock(clock), .in1(R7765));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7944 (.out1(R7945), .clock(clock), .in1(R7944));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8118 (.out1(R8119), .clock(clock), .in1(R8118));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8339 (.out1(R8340), .clock(clock), .in1(R8339));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8505 (.out1(R8506), .clock(clock), .in1(R8505));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8666 (.out1(R8667), .clock(clock), .in1(R8666));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8874 (.out1(R8875), .clock(clock), .in1(R8874));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9027 (.out1(R9028), .clock(clock), .in1(R9027));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9175 (.out1(R9176), .clock(clock), .in1(R9175));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9368 (.out1(R9369), .clock(clock), .in1(_767));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9369 (.out1(R9370), .clock(clock), .in1(_686));
  SRAM op712 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_687),.ADR(R9370));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op793 (.out1(_768), .in1(R9369), .in2(6 'd 56));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3793 (.out1(R3794), .clock(clock), .in1(R3793));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4049 (.out1(R4050), .clock(clock), .in1(R4049));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4304 (.out1(R4305), .clock(clock), .in1(R4304));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4549 (.out1(R4550), .clock(clock), .in1(R4549));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4789 (.out1(R4790), .clock(clock), .in1(R4789));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5076 (.out1(R5077), .clock(clock), .in1(R5076));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5308 (.out1(R5309), .clock(clock), .in1(R5308));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5535 (.out1(R5536), .clock(clock), .in1(R5535));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5809 (.out1(R5810), .clock(clock), .in1(R5809));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6027 (.out1(R6028), .clock(clock), .in1(R6027));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6240 (.out1(R6241), .clock(clock), .in1(R6240));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6501 (.out1(R6502), .clock(clock), .in1(R6501));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6706 (.out1(R6707), .clock(clock), .in1(R6706));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6906 (.out1(R6907), .clock(clock), .in1(R6906));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7153 (.out1(R7154), .clock(clock), .in1(R7153));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7345 (.out1(R7346), .clock(clock), .in1(R7345));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7532 (.out1(R7533), .clock(clock), .in1(R7532));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7766 (.out1(R7767), .clock(clock), .in1(R7766));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7945 (.out1(R7946), .clock(clock), .in1(R7945));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8119 (.out1(R8120), .clock(clock), .in1(R8119));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8340 (.out1(R8341), .clock(clock), .in1(R8340));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8506 (.out1(R8507), .clock(clock), .in1(R8506));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8667 (.out1(R8668), .clock(clock), .in1(R8667));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8875 (.out1(R8876), .clock(clock), .in1(R8875));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9028 (.out1(R9029), .clock(clock), .in1(R9028));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9176 (.out1(R9177), .clock(clock), .in1(R9176));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9370 (.out1(R9371), .clock(clock), .in1(_687));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9371 (.out1(R9372), .clock(clock), .in1(_768));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op794 (.out1(_769), .in1(R9372));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op795 (.out1(_770), .in1(R9371), .in2(_769));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op796 (.out1(idx_3601), .in1(_770), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3794 (.out1(R3795), .clock(clock), .in1(R3794));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4050 (.out1(R4051), .clock(clock), .in1(R4050));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4305 (.out1(R4306), .clock(clock), .in1(R4305));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4550 (.out1(R4551), .clock(clock), .in1(R4550));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4790 (.out1(R4791), .clock(clock), .in1(R4790));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5077 (.out1(R5078), .clock(clock), .in1(R5077));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5309 (.out1(R5310), .clock(clock), .in1(R5309));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5536 (.out1(R5537), .clock(clock), .in1(R5536));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5810 (.out1(R5811), .clock(clock), .in1(R5810));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6028 (.out1(R6029), .clock(clock), .in1(R6028));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6241 (.out1(R6242), .clock(clock), .in1(R6241));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6502 (.out1(R6503), .clock(clock), .in1(R6502));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6707 (.out1(R6708), .clock(clock), .in1(R6707));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6907 (.out1(R6908), .clock(clock), .in1(R6907));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7154 (.out1(R7155), .clock(clock), .in1(R7154));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7346 (.out1(R7347), .clock(clock), .in1(R7346));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7533 (.out1(R7534), .clock(clock), .in1(R7533));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7767 (.out1(R7768), .clock(clock), .in1(R7767));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7946 (.out1(R7947), .clock(clock), .in1(R7946));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8120 (.out1(R8121), .clock(clock), .in1(R8120));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8341 (.out1(R8342), .clock(clock), .in1(R8341));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8507 (.out1(R8508), .clock(clock), .in1(R8507));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8668 (.out1(R8669), .clock(clock), .in1(R8668));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8876 (.out1(R8877), .clock(clock), .in1(R8876));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9029 (.out1(R9030), .clock(clock), .in1(R9029));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9177 (.out1(R9178), .clock(clock), .in1(R9177));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9372 (.out1(R9373), .clock(clock), .in1(idx_3601));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op799 (.out1(_772), .in1(R9373));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op800 (.out1(_773), .in1(_772), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3795 (.out1(R3796), .clock(clock), .in1(R3795));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4051 (.out1(R4052), .clock(clock), .in1(R4051));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4306 (.out1(R4307), .clock(clock), .in1(R4306));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4551 (.out1(R4552), .clock(clock), .in1(R4551));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4791 (.out1(R4792), .clock(clock), .in1(R4791));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5078 (.out1(R5079), .clock(clock), .in1(R5078));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5310 (.out1(R5311), .clock(clock), .in1(R5310));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5537 (.out1(R5538), .clock(clock), .in1(R5537));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5811 (.out1(R5812), .clock(clock), .in1(R5811));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6029 (.out1(R6030), .clock(clock), .in1(R6029));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6242 (.out1(R6243), .clock(clock), .in1(R6242));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6503 (.out1(R6504), .clock(clock), .in1(R6503));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6708 (.out1(R6709), .clock(clock), .in1(R6708));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6908 (.out1(R6909), .clock(clock), .in1(R6908));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7155 (.out1(R7156), .clock(clock), .in1(R7155));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7347 (.out1(R7348), .clock(clock), .in1(R7347));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7534 (.out1(R7535), .clock(clock), .in1(R7534));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7768 (.out1(R7769), .clock(clock), .in1(R7768));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7947 (.out1(R7948), .clock(clock), .in1(R7947));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8121 (.out1(R8122), .clock(clock), .in1(R8121));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8342 (.out1(R8343), .clock(clock), .in1(R8342));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8508 (.out1(R8509), .clock(clock), .in1(R8508));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8669 (.out1(R8670), .clock(clock), .in1(R8669));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8877 (.out1(R8878), .clock(clock), .in1(R8877));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9030 (.out1(R9031), .clock(clock), .in1(R9030));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9178 (.out1(R9179), .clock(clock), .in1(R9178));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9373 (.out1(R9374), .clock(clock), .in1(R9373));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9513 (.out1(R9514), .clock(clock), .in1(_773));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op801 (.out1(_774), .in1(vec64_3604_D), .in2(R9514));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3796 (.out1(R3797), .clock(clock), .in1(R3796));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4052 (.out1(R4053), .clock(clock), .in1(R4052));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4307 (.out1(R4308), .clock(clock), .in1(R4307));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4552 (.out1(R4553), .clock(clock), .in1(R4552));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4792 (.out1(R4793), .clock(clock), .in1(R4792));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5079 (.out1(R5080), .clock(clock), .in1(R5079));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5311 (.out1(R5312), .clock(clock), .in1(R5311));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5538 (.out1(R5539), .clock(clock), .in1(R5538));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5812 (.out1(R5813), .clock(clock), .in1(R5812));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6030 (.out1(R6031), .clock(clock), .in1(R6030));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6243 (.out1(R6244), .clock(clock), .in1(R6243));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6504 (.out1(R6505), .clock(clock), .in1(R6504));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6709 (.out1(R6710), .clock(clock), .in1(R6709));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6909 (.out1(R6910), .clock(clock), .in1(R6909));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7156 (.out1(R7157), .clock(clock), .in1(R7156));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7348 (.out1(R7349), .clock(clock), .in1(R7348));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7535 (.out1(R7536), .clock(clock), .in1(R7535));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7769 (.out1(R7770), .clock(clock), .in1(R7769));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7948 (.out1(R7949), .clock(clock), .in1(R7948));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8122 (.out1(R8123), .clock(clock), .in1(R8122));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8343 (.out1(R8344), .clock(clock), .in1(R8343));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8509 (.out1(R8510), .clock(clock), .in1(R8509));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8670 (.out1(R8671), .clock(clock), .in1(R8670));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8878 (.out1(R8879), .clock(clock), .in1(R8878));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9031 (.out1(R9032), .clock(clock), .in1(R9031));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9179 (.out1(R9180), .clock(clock), .in1(R9179));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9374 (.out1(R9375), .clock(clock), .in1(R9374));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9514 (.out1(R9515), .clock(clock), .in1(_774));
  SRAM op802 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_775),.ADR(R9515));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3797 (.out1(R3798), .clock(clock), .in1(R3797));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4053 (.out1(R4054), .clock(clock), .in1(R4053));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4308 (.out1(R4309), .clock(clock), .in1(R4308));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4553 (.out1(R4554), .clock(clock), .in1(R4553));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4793 (.out1(R4794), .clock(clock), .in1(R4793));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5080 (.out1(R5081), .clock(clock), .in1(R5080));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5312 (.out1(R5313), .clock(clock), .in1(R5312));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5539 (.out1(R5540), .clock(clock), .in1(R5539));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5813 (.out1(R5814), .clock(clock), .in1(R5813));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6031 (.out1(R6032), .clock(clock), .in1(R6031));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6244 (.out1(R6245), .clock(clock), .in1(R6244));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6505 (.out1(R6506), .clock(clock), .in1(R6505));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6710 (.out1(R6711), .clock(clock), .in1(R6710));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6910 (.out1(R6911), .clock(clock), .in1(R6910));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7157 (.out1(R7158), .clock(clock), .in1(R7157));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7349 (.out1(R7350), .clock(clock), .in1(R7349));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7536 (.out1(R7537), .clock(clock), .in1(R7536));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7770 (.out1(R7771), .clock(clock), .in1(R7770));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7949 (.out1(R7950), .clock(clock), .in1(R7949));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8123 (.out1(R8124), .clock(clock), .in1(R8123));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8344 (.out1(R8345), .clock(clock), .in1(R8344));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8510 (.out1(R8511), .clock(clock), .in1(R8510));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8671 (.out1(R8672), .clock(clock), .in1(R8671));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8879 (.out1(R8880), .clock(clock), .in1(R8879));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9032 (.out1(R9033), .clock(clock), .in1(R9032));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9180 (.out1(R9181), .clock(clock), .in1(R9180));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9375 (.out1(R9376), .clock(clock), .in1(R9375));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9515 (.out1(R9516), .clock(clock), .in1(_775));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op797 (.out1(_771), .in1(ip2_3602_D), .in2(6 'd 58));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op798 (.out1(off_3603), .in1(_771));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op803 (.out1(_776), .in1(R9516), .in2(off_3603));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3798 (.out1(R3799), .clock(clock), .in1(R3798));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4054 (.out1(R4055), .clock(clock), .in1(R4054));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4309 (.out1(R4310), .clock(clock), .in1(R4309));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4554 (.out1(R4555), .clock(clock), .in1(R4554));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4794 (.out1(R4795), .clock(clock), .in1(R4794));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5081 (.out1(R5082), .clock(clock), .in1(R5081));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5313 (.out1(R5314), .clock(clock), .in1(R5313));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5540 (.out1(R5541), .clock(clock), .in1(R5540));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5814 (.out1(R5815), .clock(clock), .in1(R5814));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6032 (.out1(R6033), .clock(clock), .in1(R6032));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6245 (.out1(R6246), .clock(clock), .in1(R6245));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6506 (.out1(R6507), .clock(clock), .in1(R6506));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6711 (.out1(R6712), .clock(clock), .in1(R6711));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6911 (.out1(R6912), .clock(clock), .in1(R6911));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7158 (.out1(R7159), .clock(clock), .in1(R7158));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7350 (.out1(R7351), .clock(clock), .in1(R7350));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7537 (.out1(R7538), .clock(clock), .in1(R7537));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7771 (.out1(R7772), .clock(clock), .in1(R7771));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7950 (.out1(R7951), .clock(clock), .in1(R7950));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8124 (.out1(R8125), .clock(clock), .in1(R8124));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8345 (.out1(R8346), .clock(clock), .in1(R8345));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8511 (.out1(R8512), .clock(clock), .in1(R8511));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8672 (.out1(R8673), .clock(clock), .in1(R8672));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8880 (.out1(R8881), .clock(clock), .in1(R8880));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9033 (.out1(R9034), .clock(clock), .in1(R9033));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9181 (.out1(R9182), .clock(clock), .in1(R9181));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9376 (.out1(R9377), .clock(clock), .in1(R9376));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9516 (.out1(R9517), .clock(clock), .in1(off_3603));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9651 (.out1(R9652), .clock(clock), .in1(_776));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op804 (.out1(_777), .in1(R9652), .in2(1 'd 1));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op805 (.out1(ifout805), .in1(_777), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op873 (.out1(_845), .in1(R9377));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op866 (.out1(_838), .in1(R9377));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op855 (.out1(_827), .in1(R9377));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op835 (.out1(_807), .in1(R9377));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op874 (.out1(_846), .in1(_845), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op867 (.out1(_839), .in1(_838), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op856 (.out1(_828), .in1(_827), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op836 (.out1(_808), .in1(_807), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3799 (.out1(R3800), .clock(clock), .in1(R3799));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4055 (.out1(R4056), .clock(clock), .in1(R4055));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4310 (.out1(R4311), .clock(clock), .in1(R4310));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4555 (.out1(R4556), .clock(clock), .in1(R4555));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4795 (.out1(R4796), .clock(clock), .in1(R4795));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5082 (.out1(R5083), .clock(clock), .in1(R5082));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5314 (.out1(R5315), .clock(clock), .in1(R5314));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5541 (.out1(R5542), .clock(clock), .in1(R5541));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5815 (.out1(R5816), .clock(clock), .in1(R5815));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6033 (.out1(R6034), .clock(clock), .in1(R6033));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6246 (.out1(R6247), .clock(clock), .in1(R6246));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6507 (.out1(R6508), .clock(clock), .in1(R6507));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6712 (.out1(R6713), .clock(clock), .in1(R6712));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6912 (.out1(R6913), .clock(clock), .in1(R6912));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7159 (.out1(R7160), .clock(clock), .in1(R7159));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7351 (.out1(R7352), .clock(clock), .in1(R7351));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7538 (.out1(R7539), .clock(clock), .in1(R7538));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7772 (.out1(R7773), .clock(clock), .in1(R7772));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7951 (.out1(R7952), .clock(clock), .in1(R7951));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8125 (.out1(R8126), .clock(clock), .in1(R8125));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8346 (.out1(R8347), .clock(clock), .in1(R8346));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8512 (.out1(R8513), .clock(clock), .in1(R8512));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8673 (.out1(R8674), .clock(clock), .in1(R8673));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8881 (.out1(R8882), .clock(clock), .in1(R8881));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9034 (.out1(R9035), .clock(clock), .in1(R9034));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9182 (.out1(R9183), .clock(clock), .in1(R9182));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9377 (.out1(R9378), .clock(clock), .in1(R9377));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9517 (.out1(R9518), .clock(clock), .in1(R9517));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9652 (.out1(R9653), .clock(clock), .in1(ifout805));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9794 (.out1(R9795), .clock(clock), .in1(_846));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9795 (.out1(R9796), .clock(clock), .in1(_839));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9796 (.out1(R9797), .clock(clock), .in1(_828));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9797 (.out1(R9798), .clock(clock), .in1(_808));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op848 (.out1(_820), .in1(R9378));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op828 (.out1(_800), .in1(R9378));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op817 (.out1(_789), .in1(R9378));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op810 (.out1(_782), .in1(R9378));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op877 (.out1(_849), .in1(2 'd 2), .in2(R9518));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op849 (.out1(_821), .in1(_820), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op829 (.out1(_801), .in1(_800), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op818 (.out1(_790), .in1(_789), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op811 (.out1(_783), .in1(_782), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op875 (.out1(_847), .in1(vec64_3604_D), .in2(R9795));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op868 (.out1(_840), .in1(vec64_3604_D), .in2(R9796));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op857 (.out1(_829), .in1(vec64_3604_D), .in2(R9797));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op837 (.out1(_809), .in1(vec64_3604_D), .in2(R9798));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3800 (.out1(R3801), .clock(clock), .in1(R3800));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4056 (.out1(R4057), .clock(clock), .in1(R4056));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4311 (.out1(R4312), .clock(clock), .in1(R4311));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4556 (.out1(R4557), .clock(clock), .in1(R4556));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4796 (.out1(R4797), .clock(clock), .in1(R4796));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5083 (.out1(R5084), .clock(clock), .in1(R5083));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5315 (.out1(R5316), .clock(clock), .in1(R5315));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5542 (.out1(R5543), .clock(clock), .in1(R5542));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5816 (.out1(R5817), .clock(clock), .in1(R5816));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6034 (.out1(R6035), .clock(clock), .in1(R6034));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6247 (.out1(R6248), .clock(clock), .in1(R6247));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6508 (.out1(R6509), .clock(clock), .in1(R6508));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6713 (.out1(R6714), .clock(clock), .in1(R6713));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6913 (.out1(R6914), .clock(clock), .in1(R6913));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7160 (.out1(R7161), .clock(clock), .in1(R7160));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7352 (.out1(R7353), .clock(clock), .in1(R7352));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7539 (.out1(R7540), .clock(clock), .in1(R7539));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7773 (.out1(R7774), .clock(clock), .in1(R7773));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7952 (.out1(R7953), .clock(clock), .in1(R7952));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8126 (.out1(R8127), .clock(clock), .in1(R8126));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8347 (.out1(R8348), .clock(clock), .in1(R8347));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8513 (.out1(R8514), .clock(clock), .in1(R8513));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8674 (.out1(R8675), .clock(clock), .in1(R8674));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8882 (.out1(R8883), .clock(clock), .in1(R8882));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9035 (.out1(R9036), .clock(clock), .in1(R9035));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9183 (.out1(R9184), .clock(clock), .in1(R9183));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9378 (.out1(R9379), .clock(clock), .in1(R9378));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9518 (.out1(R9519), .clock(clock), .in1(R9518));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9653 (.out1(R9654), .clock(clock), .in1(R9653));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9798 (.out1(R9799), .clock(clock), .in1(_849));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9799 (.out1(R9800), .clock(clock), .in1(_821));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9800 (.out1(R9801), .clock(clock), .in1(_801));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9801 (.out1(R9802), .clock(clock), .in1(_790));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9802 (.out1(R9803), .clock(clock), .in1(_783));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9803 (.out1(R9804), .clock(clock), .in1(_847));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9804 (.out1(R9805), .clock(clock), .in1(_840));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9805 (.out1(R9806), .clock(clock), .in1(_829));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9806 (.out1(R9807), .clock(clock), .in1(_809));
  SRAM op876 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_848),.ADR(R9804));
  SRAM op869 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_841),.ADR(R9805));
  SRAM op858 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_830),.ADR(R9806));
  SRAM op838 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_810),.ADR(R9807));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op870 (.out1(_842), .in1(2 'd 2), .in2(R9519));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op859 (.out1(_831), .in1(2 'd 2), .in2(R9519));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op852 (.out1(_824), .in1(2 'd 2), .in2(R9519));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op839 (.out1(_811), .in1(2 'd 2), .in2(R9519));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op832 (.out1(_804), .in1(2 'd 2), .in2(R9519));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op821 (.out1(_793), .in1(2 'd 2), .in2(R9519));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op850 (.out1(_822), .in1(vec64_3604_D), .in2(R9800));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op830 (.out1(_802), .in1(vec64_3604_D), .in2(R9801));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op819 (.out1(_791), .in1(vec64_3604_D), .in2(R9802));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op812 (.out1(_784), .in1(vec64_3604_D), .in2(R9803));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op878 (.out1(_850), .in1(R9799), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3801 (.out1(R3802), .clock(clock), .in1(R3801));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4057 (.out1(R4058), .clock(clock), .in1(R4057));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4312 (.out1(R4313), .clock(clock), .in1(R4312));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4557 (.out1(R4558), .clock(clock), .in1(R4557));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4797 (.out1(R4798), .clock(clock), .in1(R4797));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5084 (.out1(R5085), .clock(clock), .in1(R5084));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5316 (.out1(R5317), .clock(clock), .in1(R5316));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5543 (.out1(R5544), .clock(clock), .in1(R5543));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5817 (.out1(R5818), .clock(clock), .in1(R5817));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6035 (.out1(R6036), .clock(clock), .in1(R6035));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6248 (.out1(R6249), .clock(clock), .in1(R6248));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6509 (.out1(R6510), .clock(clock), .in1(R6509));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6714 (.out1(R6715), .clock(clock), .in1(R6714));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6914 (.out1(R6915), .clock(clock), .in1(R6914));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7161 (.out1(R7162), .clock(clock), .in1(R7161));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7353 (.out1(R7354), .clock(clock), .in1(R7353));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7540 (.out1(R7541), .clock(clock), .in1(R7540));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7774 (.out1(R7775), .clock(clock), .in1(R7774));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7953 (.out1(R7954), .clock(clock), .in1(R7953));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8127 (.out1(R8128), .clock(clock), .in1(R8127));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8348 (.out1(R8349), .clock(clock), .in1(R8348));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8514 (.out1(R8515), .clock(clock), .in1(R8514));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8675 (.out1(R8676), .clock(clock), .in1(R8675));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8883 (.out1(R8884), .clock(clock), .in1(R8883));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9036 (.out1(R9037), .clock(clock), .in1(R9036));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9184 (.out1(R9185), .clock(clock), .in1(R9184));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9379 (.out1(R9380), .clock(clock), .in1(R9379));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9519 (.out1(R9520), .clock(clock), .in1(R9519));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9654 (.out1(R9655), .clock(clock), .in1(R9654));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9807 (.out1(R9808), .clock(clock), .in1(_848));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9808 (.out1(R9809), .clock(clock), .in1(_841));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9809 (.out1(R9810), .clock(clock), .in1(_830));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9810 (.out1(R9811), .clock(clock), .in1(_810));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9811 (.out1(R9812), .clock(clock), .in1(_842));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9812 (.out1(R9813), .clock(clock), .in1(_831));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9813 (.out1(R9814), .clock(clock), .in1(_824));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9814 (.out1(R9815), .clock(clock), .in1(_811));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9815 (.out1(R9816), .clock(clock), .in1(_804));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9816 (.out1(R9817), .clock(clock), .in1(_793));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9817 (.out1(R9818), .clock(clock), .in1(_822));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9818 (.out1(R9819), .clock(clock), .in1(_802));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9819 (.out1(R9820), .clock(clock), .in1(_791));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9820 (.out1(R9821), .clock(clock), .in1(_784));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9821 (.out1(R9822), .clock(clock), .in1(_850));
  SRAM op851 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_823),.ADR(R9818));
  SRAM op831 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_803),.ADR(R9819));
  SRAM op820 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_792),.ADR(R9820));
  SRAM op813 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_785),.ADR(R9821));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op879 (.out1(_851), .in1(R9808), .in2(R9822));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op880 (.out1(_852), .in1(_851), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op871 (.out1(_843), .in1(R9812), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op860 (.out1(_832), .in1(R9813), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op840 (.out1(_812), .in1(R9815), .in2(64 'd 18446744073709551615));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op814 (.out1(_786), .in1(2 'd 2), .in2(R9520));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op881 (.out1(_853), .in1(_852), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op872 (.out1(_844), .in1(R9809), .in2(_843));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op861 (.out1(_833), .in1(R9810), .in2(_832));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op841 (.out1(_813), .in1(R9811), .in2(_812));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op882 (.out1(_854), .in1(_844), .in2(_853));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op862 (.out1(_834), .in1(_833), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op853 (.out1(_825), .in1(R9814), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op842 (.out1(_814), .in1(_813), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op833 (.out1(_805), .in1(R9816), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op822 (.out1(_794), .in1(R9817), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3802 (.out1(R3803), .clock(clock), .in1(R3802));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4058 (.out1(R4059), .clock(clock), .in1(R4058));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4313 (.out1(R4314), .clock(clock), .in1(R4313));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4558 (.out1(R4559), .clock(clock), .in1(R4558));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4798 (.out1(R4799), .clock(clock), .in1(R4798));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5085 (.out1(R5086), .clock(clock), .in1(R5085));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5317 (.out1(R5318), .clock(clock), .in1(R5317));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5544 (.out1(R5545), .clock(clock), .in1(R5544));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5818 (.out1(R5819), .clock(clock), .in1(R5818));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6036 (.out1(R6037), .clock(clock), .in1(R6036));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6249 (.out1(R6250), .clock(clock), .in1(R6249));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6510 (.out1(R6511), .clock(clock), .in1(R6510));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6715 (.out1(R6716), .clock(clock), .in1(R6715));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6915 (.out1(R6916), .clock(clock), .in1(R6915));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7162 (.out1(R7163), .clock(clock), .in1(R7162));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7354 (.out1(R7355), .clock(clock), .in1(R7354));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7541 (.out1(R7542), .clock(clock), .in1(R7541));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7775 (.out1(R7776), .clock(clock), .in1(R7775));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7954 (.out1(R7955), .clock(clock), .in1(R7954));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8128 (.out1(R8129), .clock(clock), .in1(R8128));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8349 (.out1(R8350), .clock(clock), .in1(R8349));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8515 (.out1(R8516), .clock(clock), .in1(R8515));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8676 (.out1(R8677), .clock(clock), .in1(R8676));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8884 (.out1(R8885), .clock(clock), .in1(R8884));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9037 (.out1(R9038), .clock(clock), .in1(R9037));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9185 (.out1(R9186), .clock(clock), .in1(R9185));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9380 (.out1(R9381), .clock(clock), .in1(R9380));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9520 (.out1(R9521), .clock(clock), .in1(R9520));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9655 (.out1(R9656), .clock(clock), .in1(R9655));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9822 (.out1(R9823), .clock(clock), .in1(_823));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9823 (.out1(R9824), .clock(clock), .in1(_803));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9824 (.out1(R9825), .clock(clock), .in1(_792));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9825 (.out1(R9826), .clock(clock), .in1(_785));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9826 (.out1(R9827), .clock(clock), .in1(_786));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9827 (.out1(R9828), .clock(clock), .in1(_854));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9828 (.out1(R9829), .clock(clock), .in1(_834));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9829 (.out1(R9830), .clock(clock), .in1(_825));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9830 (.out1(R9831), .clock(clock), .in1(_814));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9831 (.out1(R9832), .clock(clock), .in1(_805));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9832 (.out1(R9833), .clock(clock), .in1(_794));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op863 (.out1(_835), .in1(R9829), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op854 (.out1(_826), .in1(R9823), .in2(R9830));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op823 (.out1(_795), .in1(R9825), .in2(R9833));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op883 (.out1(_855), .in1(R9828), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op864 (.out1(_836), .in1(_826), .in2(_835));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op843 (.out1(_815), .in1(R9831), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op834 (.out1(_806), .in1(R9824), .in2(R9832));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op824 (.out1(_796), .in1(_795), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op815 (.out1(_787), .in1(R9827), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op844 (.out1(_816), .in1(_806), .in2(_815));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op884 (.out1(_856), .in1(_855), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op865 (.out1(_837), .in1(_836), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op825 (.out1(_797), .in1(_796), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op816 (.out1(_788), .in1(R9826), .in2(_787));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op885 (.out1(_857), .in1(_837), .in2(_856));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op845 (.out1(_817), .in1(_816), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op826 (.out1(_798), .in1(_788), .in2(_797));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3803 (.out1(R3804), .clock(clock), .in1(R3803));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4059 (.out1(R4060), .clock(clock), .in1(R4059));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4314 (.out1(R4315), .clock(clock), .in1(R4314));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4559 (.out1(R4560), .clock(clock), .in1(R4559));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4799 (.out1(R4800), .clock(clock), .in1(R4799));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5086 (.out1(R5087), .clock(clock), .in1(R5086));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5318 (.out1(R5319), .clock(clock), .in1(R5318));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5545 (.out1(R5546), .clock(clock), .in1(R5545));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5819 (.out1(R5820), .clock(clock), .in1(R5819));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6037 (.out1(R6038), .clock(clock), .in1(R6037));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6250 (.out1(R6251), .clock(clock), .in1(R6250));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6511 (.out1(R6512), .clock(clock), .in1(R6511));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6716 (.out1(R6717), .clock(clock), .in1(R6716));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6916 (.out1(R6917), .clock(clock), .in1(R6916));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7163 (.out1(R7164), .clock(clock), .in1(R7163));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7355 (.out1(R7356), .clock(clock), .in1(R7355));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7542 (.out1(R7543), .clock(clock), .in1(R7542));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7776 (.out1(R7777), .clock(clock), .in1(R7776));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7955 (.out1(R7956), .clock(clock), .in1(R7955));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8129 (.out1(R8130), .clock(clock), .in1(R8129));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8350 (.out1(R8351), .clock(clock), .in1(R8350));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8516 (.out1(R8517), .clock(clock), .in1(R8516));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8677 (.out1(R8678), .clock(clock), .in1(R8677));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8885 (.out1(R8886), .clock(clock), .in1(R8885));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9038 (.out1(R9039), .clock(clock), .in1(R9038));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9186 (.out1(R9187), .clock(clock), .in1(R9186));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9381 (.out1(R9382), .clock(clock), .in1(R9381));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9521 (.out1(R9522), .clock(clock), .in1(R9521));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9656 (.out1(R9657), .clock(clock), .in1(R9656));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9833 (.out1(R9834), .clock(clock), .in1(_857));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9834 (.out1(R9835), .clock(clock), .in1(_817));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9835 (.out1(R9836), .clock(clock), .in1(_798));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op806 (.out1(_778), .in1(R9382));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op846 (.out1(_818), .in1(R9835), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op827 (.out1(_799), .in1(R9836), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op886 (.out1(_858), .in1(R9834), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op847 (.out1(_819), .in1(_799), .in2(_818));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op807 (.out1(_779), .in1(_778), .in2(2 'd 2));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op887 (.out1(_859), .in1(_819), .in2(_858));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op888 (.out1(_860), .in1(_859), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3804 (.out1(R3805), .clock(clock), .in1(R3804));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4060 (.out1(R4061), .clock(clock), .in1(R4060));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4315 (.out1(R4316), .clock(clock), .in1(R4315));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4560 (.out1(R4561), .clock(clock), .in1(R4560));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4800 (.out1(R4801), .clock(clock), .in1(R4800));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5087 (.out1(R5088), .clock(clock), .in1(R5087));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5319 (.out1(R5320), .clock(clock), .in1(R5319));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5546 (.out1(R5547), .clock(clock), .in1(R5546));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5820 (.out1(R5821), .clock(clock), .in1(R5820));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6038 (.out1(R6039), .clock(clock), .in1(R6038));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6251 (.out1(R6252), .clock(clock), .in1(R6251));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6512 (.out1(R6513), .clock(clock), .in1(R6512));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6717 (.out1(R6718), .clock(clock), .in1(R6717));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6917 (.out1(R6918), .clock(clock), .in1(R6917));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7164 (.out1(R7165), .clock(clock), .in1(R7164));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7356 (.out1(R7357), .clock(clock), .in1(R7356));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7543 (.out1(R7544), .clock(clock), .in1(R7543));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7777 (.out1(R7778), .clock(clock), .in1(R7777));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7956 (.out1(R7957), .clock(clock), .in1(R7956));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8130 (.out1(R8131), .clock(clock), .in1(R8130));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8351 (.out1(R8352), .clock(clock), .in1(R8351));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8517 (.out1(R8518), .clock(clock), .in1(R8517));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8678 (.out1(R8679), .clock(clock), .in1(R8678));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8886 (.out1(R8887), .clock(clock), .in1(R8886));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9039 (.out1(R9040), .clock(clock), .in1(R9039));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9187 (.out1(R9188), .clock(clock), .in1(R9187));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9382 (.out1(R9383), .clock(clock), .in1(R9382));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9522 (.out1(R9523), .clock(clock), .in1(R9522));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9657 (.out1(R9658), .clock(clock), .in1(R9657));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9836 (.out1(R9837), .clock(clock), .in1(_779));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9837 (.out1(R9838), .clock(clock), .in1(_860));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op889 (.out1(_861), .in1(R9838), .in2(57 'd 72340172838076673));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op808 (.out1(_780), .in1(base0_64_3609_D), .in2(R9837));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3805 (.out1(R3806), .clock(clock), .in1(R3805));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4061 (.out1(R4062), .clock(clock), .in1(R4061));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4316 (.out1(R4317), .clock(clock), .in1(R4316));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4561 (.out1(R4562), .clock(clock), .in1(R4561));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4801 (.out1(R4802), .clock(clock), .in1(R4801));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5088 (.out1(R5089), .clock(clock), .in1(R5088));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5320 (.out1(R5321), .clock(clock), .in1(R5320));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5547 (.out1(R5548), .clock(clock), .in1(R5547));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5821 (.out1(R5822), .clock(clock), .in1(R5821));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6039 (.out1(R6040), .clock(clock), .in1(R6039));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6252 (.out1(R6253), .clock(clock), .in1(R6252));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6513 (.out1(R6514), .clock(clock), .in1(R6513));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6718 (.out1(R6719), .clock(clock), .in1(R6718));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6918 (.out1(R6919), .clock(clock), .in1(R6918));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7165 (.out1(R7166), .clock(clock), .in1(R7165));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7357 (.out1(R7358), .clock(clock), .in1(R7357));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7544 (.out1(R7545), .clock(clock), .in1(R7544));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7778 (.out1(R7779), .clock(clock), .in1(R7778));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7957 (.out1(R7958), .clock(clock), .in1(R7957));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8131 (.out1(R8132), .clock(clock), .in1(R8131));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8352 (.out1(R8353), .clock(clock), .in1(R8352));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8518 (.out1(R8519), .clock(clock), .in1(R8518));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8679 (.out1(R8680), .clock(clock), .in1(R8679));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8887 (.out1(R8888), .clock(clock), .in1(R8887));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9040 (.out1(R9041), .clock(clock), .in1(R9040));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9188 (.out1(R9189), .clock(clock), .in1(R9188));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9383 (.out1(R9384), .clock(clock), .in1(R9383));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9523 (.out1(R9524), .clock(clock), .in1(R9523));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9658 (.out1(R9659), .clock(clock), .in1(R9658));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9838 (.out1(R9839), .clock(clock), .in1(_861));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9839 (.out1(R9840), .clock(clock), .in1(_780));
  SRAM op809 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_781),.ADR(R9840));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op890 (.out1(_862), .in1(R9839), .in2(6 'd 56));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3806 (.out1(R3807), .clock(clock), .in1(R3806));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4062 (.out1(R4063), .clock(clock), .in1(R4062));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4317 (.out1(R4318), .clock(clock), .in1(R4317));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4562 (.out1(R4563), .clock(clock), .in1(R4562));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4802 (.out1(R4803), .clock(clock), .in1(R4802));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5089 (.out1(R5090), .clock(clock), .in1(R5089));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5321 (.out1(R5322), .clock(clock), .in1(R5321));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5548 (.out1(R5549), .clock(clock), .in1(R5548));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5822 (.out1(R5823), .clock(clock), .in1(R5822));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6040 (.out1(R6041), .clock(clock), .in1(R6040));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6253 (.out1(R6254), .clock(clock), .in1(R6253));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6514 (.out1(R6515), .clock(clock), .in1(R6514));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6719 (.out1(R6720), .clock(clock), .in1(R6719));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6919 (.out1(R6920), .clock(clock), .in1(R6919));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7166 (.out1(R7167), .clock(clock), .in1(R7166));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7358 (.out1(R7359), .clock(clock), .in1(R7358));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7545 (.out1(R7546), .clock(clock), .in1(R7545));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7779 (.out1(R7780), .clock(clock), .in1(R7779));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7958 (.out1(R7959), .clock(clock), .in1(R7958));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8132 (.out1(R8133), .clock(clock), .in1(R8132));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8353 (.out1(R8354), .clock(clock), .in1(R8353));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8519 (.out1(R8520), .clock(clock), .in1(R8519));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8680 (.out1(R8681), .clock(clock), .in1(R8680));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8888 (.out1(R8889), .clock(clock), .in1(R8888));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9041 (.out1(R9042), .clock(clock), .in1(R9041));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9189 (.out1(R9190), .clock(clock), .in1(R9189));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9384 (.out1(R9385), .clock(clock), .in1(R9384));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9524 (.out1(R9525), .clock(clock), .in1(R9524));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9659 (.out1(R9660), .clock(clock), .in1(R9659));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9840 (.out1(R9841), .clock(clock), .in1(_781));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9841 (.out1(R9842), .clock(clock), .in1(_862));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op891 (.out1(_863), .in1(R9842));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op892 (.out1(_864), .in1(R9841), .in2(_863));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op893 (.out1(idx_3610), .in1(_864), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3807 (.out1(R3808), .clock(clock), .in1(R3807));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4063 (.out1(R4064), .clock(clock), .in1(R4063));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4318 (.out1(R4319), .clock(clock), .in1(R4318));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4563 (.out1(R4564), .clock(clock), .in1(R4563));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4803 (.out1(R4804), .clock(clock), .in1(R4803));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5090 (.out1(R5091), .clock(clock), .in1(R5090));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5322 (.out1(R5323), .clock(clock), .in1(R5322));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5549 (.out1(R5550), .clock(clock), .in1(R5549));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5823 (.out1(R5824), .clock(clock), .in1(R5823));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6041 (.out1(R6042), .clock(clock), .in1(R6041));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6254 (.out1(R6255), .clock(clock), .in1(R6254));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6515 (.out1(R6516), .clock(clock), .in1(R6515));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6720 (.out1(R6721), .clock(clock), .in1(R6720));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6920 (.out1(R6921), .clock(clock), .in1(R6920));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7167 (.out1(R7168), .clock(clock), .in1(R7167));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7359 (.out1(R7360), .clock(clock), .in1(R7359));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7546 (.out1(R7547), .clock(clock), .in1(R7546));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7780 (.out1(R7781), .clock(clock), .in1(R7780));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7959 (.out1(R7960), .clock(clock), .in1(R7959));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8133 (.out1(R8134), .clock(clock), .in1(R8133));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8354 (.out1(R8355), .clock(clock), .in1(R8354));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8520 (.out1(R8521), .clock(clock), .in1(R8520));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8681 (.out1(R8682), .clock(clock), .in1(R8681));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8889 (.out1(R8890), .clock(clock), .in1(R8889));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9042 (.out1(R9043), .clock(clock), .in1(R9042));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9190 (.out1(R9191), .clock(clock), .in1(R9190));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9385 (.out1(R9386), .clock(clock), .in1(R9385));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9525 (.out1(R9526), .clock(clock), .in1(R9525));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9660 (.out1(R9661), .clock(clock), .in1(R9660));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9842 (.out1(R9843), .clock(clock), .in1(idx_3610));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op897 (.out1(_867), .in1(R9843));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op898 (.out1(_868), .in1(_867), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3808 (.out1(R3809), .clock(clock), .in1(R3808));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4064 (.out1(R4065), .clock(clock), .in1(R4064));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4319 (.out1(R4320), .clock(clock), .in1(R4319));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4564 (.out1(R4565), .clock(clock), .in1(R4564));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4804 (.out1(R4805), .clock(clock), .in1(R4804));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5091 (.out1(R5092), .clock(clock), .in1(R5091));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5323 (.out1(R5324), .clock(clock), .in1(R5323));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5550 (.out1(R5551), .clock(clock), .in1(R5550));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5824 (.out1(R5825), .clock(clock), .in1(R5824));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6042 (.out1(R6043), .clock(clock), .in1(R6042));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6255 (.out1(R6256), .clock(clock), .in1(R6255));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6516 (.out1(R6517), .clock(clock), .in1(R6516));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6721 (.out1(R6722), .clock(clock), .in1(R6721));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6921 (.out1(R6922), .clock(clock), .in1(R6921));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7168 (.out1(R7169), .clock(clock), .in1(R7168));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7360 (.out1(R7361), .clock(clock), .in1(R7360));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7547 (.out1(R7548), .clock(clock), .in1(R7547));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7781 (.out1(R7782), .clock(clock), .in1(R7781));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7960 (.out1(R7961), .clock(clock), .in1(R7960));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8134 (.out1(R8135), .clock(clock), .in1(R8134));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8355 (.out1(R8356), .clock(clock), .in1(R8355));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8521 (.out1(R8522), .clock(clock), .in1(R8521));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8682 (.out1(R8683), .clock(clock), .in1(R8682));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8890 (.out1(R8891), .clock(clock), .in1(R8890));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9043 (.out1(R9044), .clock(clock), .in1(R9043));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9191 (.out1(R9192), .clock(clock), .in1(R9191));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9386 (.out1(R9387), .clock(clock), .in1(R9386));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9526 (.out1(R9527), .clock(clock), .in1(R9526));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9661 (.out1(R9662), .clock(clock), .in1(R9661));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9843 (.out1(R9844), .clock(clock), .in1(R9843));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9970 (.out1(R9971), .clock(clock), .in1(_868));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op899 (.out1(_869), .in1(vec70_3612_D), .in2(R9971));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3809 (.out1(R3810), .clock(clock), .in1(R3809));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4065 (.out1(R4066), .clock(clock), .in1(R4065));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4320 (.out1(R4321), .clock(clock), .in1(R4320));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4565 (.out1(R4566), .clock(clock), .in1(R4565));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4805 (.out1(R4806), .clock(clock), .in1(R4805));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5092 (.out1(R5093), .clock(clock), .in1(R5092));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5324 (.out1(R5325), .clock(clock), .in1(R5324));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5551 (.out1(R5552), .clock(clock), .in1(R5551));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5825 (.out1(R5826), .clock(clock), .in1(R5825));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6043 (.out1(R6044), .clock(clock), .in1(R6043));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6256 (.out1(R6257), .clock(clock), .in1(R6256));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6517 (.out1(R6518), .clock(clock), .in1(R6517));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6722 (.out1(R6723), .clock(clock), .in1(R6722));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6922 (.out1(R6923), .clock(clock), .in1(R6922));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7169 (.out1(R7170), .clock(clock), .in1(R7169));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7361 (.out1(R7362), .clock(clock), .in1(R7361));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7548 (.out1(R7549), .clock(clock), .in1(R7548));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7782 (.out1(R7783), .clock(clock), .in1(R7782));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7961 (.out1(R7962), .clock(clock), .in1(R7961));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8135 (.out1(R8136), .clock(clock), .in1(R8135));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8356 (.out1(R8357), .clock(clock), .in1(R8356));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8522 (.out1(R8523), .clock(clock), .in1(R8522));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8683 (.out1(R8684), .clock(clock), .in1(R8683));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8891 (.out1(R8892), .clock(clock), .in1(R8891));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9044 (.out1(R9045), .clock(clock), .in1(R9044));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9192 (.out1(R9193), .clock(clock), .in1(R9192));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9387 (.out1(R9388), .clock(clock), .in1(R9387));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9527 (.out1(R9528), .clock(clock), .in1(R9527));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9662 (.out1(R9663), .clock(clock), .in1(R9662));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9844 (.out1(R9845), .clock(clock), .in1(R9844));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9971 (.out1(R9972), .clock(clock), .in1(_869));
  SRAM op900 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_870),.ADR(R9972));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3810 (.out1(R3811), .clock(clock), .in1(R3810));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4066 (.out1(R4067), .clock(clock), .in1(R4066));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4321 (.out1(R4322), .clock(clock), .in1(R4321));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4566 (.out1(R4567), .clock(clock), .in1(R4566));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4806 (.out1(R4807), .clock(clock), .in1(R4806));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5093 (.out1(R5094), .clock(clock), .in1(R5093));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5325 (.out1(R5326), .clock(clock), .in1(R5325));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5552 (.out1(R5553), .clock(clock), .in1(R5552));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5826 (.out1(R5827), .clock(clock), .in1(R5826));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6044 (.out1(R6045), .clock(clock), .in1(R6044));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6257 (.out1(R6258), .clock(clock), .in1(R6257));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6518 (.out1(R6519), .clock(clock), .in1(R6518));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6723 (.out1(R6724), .clock(clock), .in1(R6723));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6923 (.out1(R6924), .clock(clock), .in1(R6923));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7170 (.out1(R7171), .clock(clock), .in1(R7170));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7362 (.out1(R7363), .clock(clock), .in1(R7362));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7549 (.out1(R7550), .clock(clock), .in1(R7549));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7783 (.out1(R7784), .clock(clock), .in1(R7783));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7962 (.out1(R7963), .clock(clock), .in1(R7962));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8136 (.out1(R8137), .clock(clock), .in1(R8136));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8357 (.out1(R8358), .clock(clock), .in1(R8357));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8523 (.out1(R8524), .clock(clock), .in1(R8523));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8684 (.out1(R8685), .clock(clock), .in1(R8684));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8892 (.out1(R8893), .clock(clock), .in1(R8892));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9045 (.out1(R9046), .clock(clock), .in1(R9045));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9193 (.out1(R9194), .clock(clock), .in1(R9193));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9388 (.out1(R9389), .clock(clock), .in1(R9388));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9528 (.out1(R9529), .clock(clock), .in1(R9528));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9663 (.out1(R9664), .clock(clock), .in1(R9663));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9845 (.out1(R9846), .clock(clock), .in1(R9845));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op9972 (.out1(R9973), .clock(clock), .in1(_870));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op894 (.out1(_865), .in1(ip2_3602_D), .in2(6 'd 52));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op895 (.out1(_866), .in1(_865));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op896 (.out1(off_3611), .in1(_866), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op901 (.out1(_871), .in1(R9973), .in2(off_3611));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3811 (.out1(R3812), .clock(clock), .in1(R3811));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4067 (.out1(R4068), .clock(clock), .in1(R4067));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4322 (.out1(R4323), .clock(clock), .in1(R4322));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4567 (.out1(R4568), .clock(clock), .in1(R4567));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4807 (.out1(R4808), .clock(clock), .in1(R4807));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5094 (.out1(R5095), .clock(clock), .in1(R5094));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5326 (.out1(R5327), .clock(clock), .in1(R5326));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5553 (.out1(R5554), .clock(clock), .in1(R5553));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5827 (.out1(R5828), .clock(clock), .in1(R5827));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6045 (.out1(R6046), .clock(clock), .in1(R6045));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6258 (.out1(R6259), .clock(clock), .in1(R6258));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6519 (.out1(R6520), .clock(clock), .in1(R6519));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6724 (.out1(R6725), .clock(clock), .in1(R6724));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6924 (.out1(R6925), .clock(clock), .in1(R6924));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7171 (.out1(R7172), .clock(clock), .in1(R7171));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7363 (.out1(R7364), .clock(clock), .in1(R7363));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7550 (.out1(R7551), .clock(clock), .in1(R7550));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7784 (.out1(R7785), .clock(clock), .in1(R7784));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7963 (.out1(R7964), .clock(clock), .in1(R7963));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8137 (.out1(R8138), .clock(clock), .in1(R8137));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8358 (.out1(R8359), .clock(clock), .in1(R8358));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8524 (.out1(R8525), .clock(clock), .in1(R8524));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8685 (.out1(R8686), .clock(clock), .in1(R8685));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8893 (.out1(R8894), .clock(clock), .in1(R8893));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9046 (.out1(R9047), .clock(clock), .in1(R9046));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9194 (.out1(R9195), .clock(clock), .in1(R9194));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9389 (.out1(R9390), .clock(clock), .in1(R9389));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9529 (.out1(R9530), .clock(clock), .in1(R9529));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9664 (.out1(R9665), .clock(clock), .in1(R9664));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9846 (.out1(R9847), .clock(clock), .in1(R9846));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9973 (.out1(R9974), .clock(clock), .in1(off_3611));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10095 (.out1(R10096), .clock(clock), .in1(_871));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op902 (.out1(_872), .in1(R10096), .in2(1 'd 1));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op903 (.out1(ifout903), .in1(_872), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op971 (.out1(_940), .in1(R9847));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op964 (.out1(_933), .in1(R9847));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op953 (.out1(_922), .in1(R9847));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op933 (.out1(_902), .in1(R9847));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op972 (.out1(_941), .in1(_940), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op965 (.out1(_934), .in1(_933), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op954 (.out1(_923), .in1(_922), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op934 (.out1(_903), .in1(_902), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3812 (.out1(R3813), .clock(clock), .in1(R3812));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4068 (.out1(R4069), .clock(clock), .in1(R4068));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4323 (.out1(R4324), .clock(clock), .in1(R4323));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4568 (.out1(R4569), .clock(clock), .in1(R4568));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4808 (.out1(R4809), .clock(clock), .in1(R4808));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5095 (.out1(R5096), .clock(clock), .in1(R5095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5327 (.out1(R5328), .clock(clock), .in1(R5327));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5554 (.out1(R5555), .clock(clock), .in1(R5554));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5828 (.out1(R5829), .clock(clock), .in1(R5828));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6046 (.out1(R6047), .clock(clock), .in1(R6046));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6259 (.out1(R6260), .clock(clock), .in1(R6259));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6520 (.out1(R6521), .clock(clock), .in1(R6520));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6725 (.out1(R6726), .clock(clock), .in1(R6725));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6925 (.out1(R6926), .clock(clock), .in1(R6925));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7172 (.out1(R7173), .clock(clock), .in1(R7172));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7364 (.out1(R7365), .clock(clock), .in1(R7364));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7551 (.out1(R7552), .clock(clock), .in1(R7551));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7785 (.out1(R7786), .clock(clock), .in1(R7785));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7964 (.out1(R7965), .clock(clock), .in1(R7964));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8138 (.out1(R8139), .clock(clock), .in1(R8138));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8359 (.out1(R8360), .clock(clock), .in1(R8359));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8525 (.out1(R8526), .clock(clock), .in1(R8525));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8686 (.out1(R8687), .clock(clock), .in1(R8686));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8894 (.out1(R8895), .clock(clock), .in1(R8894));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9047 (.out1(R9048), .clock(clock), .in1(R9047));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9195 (.out1(R9196), .clock(clock), .in1(R9195));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9390 (.out1(R9391), .clock(clock), .in1(R9390));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9530 (.out1(R9531), .clock(clock), .in1(R9530));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9665 (.out1(R9666), .clock(clock), .in1(R9665));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9847 (.out1(R9848), .clock(clock), .in1(R9847));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9974 (.out1(R9975), .clock(clock), .in1(R9974));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10096 (.out1(R10097), .clock(clock), .in1(ifout903));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10225 (.out1(R10226), .clock(clock), .in1(_941));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10226 (.out1(R10227), .clock(clock), .in1(_934));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10227 (.out1(R10228), .clock(clock), .in1(_923));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10228 (.out1(R10229), .clock(clock), .in1(_903));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op946 (.out1(_915), .in1(R9848));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op926 (.out1(_895), .in1(R9848));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op915 (.out1(_884), .in1(R9848));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op908 (.out1(_877), .in1(R9848));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op975 (.out1(_944), .in1(2 'd 2), .in2(R9975));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op947 (.out1(_916), .in1(_915), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op927 (.out1(_896), .in1(_895), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op916 (.out1(_885), .in1(_884), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op909 (.out1(_878), .in1(_877), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op973 (.out1(_942), .in1(vec70_3612_D), .in2(R10226));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op966 (.out1(_935), .in1(vec70_3612_D), .in2(R10227));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op955 (.out1(_924), .in1(vec70_3612_D), .in2(R10228));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op935 (.out1(_904), .in1(vec70_3612_D), .in2(R10229));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3813 (.out1(R3814), .clock(clock), .in1(R3813));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4069 (.out1(R4070), .clock(clock), .in1(R4069));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4324 (.out1(R4325), .clock(clock), .in1(R4324));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4569 (.out1(R4570), .clock(clock), .in1(R4569));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4809 (.out1(R4810), .clock(clock), .in1(R4809));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5096 (.out1(R5097), .clock(clock), .in1(R5096));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5328 (.out1(R5329), .clock(clock), .in1(R5328));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5555 (.out1(R5556), .clock(clock), .in1(R5555));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5829 (.out1(R5830), .clock(clock), .in1(R5829));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6047 (.out1(R6048), .clock(clock), .in1(R6047));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6260 (.out1(R6261), .clock(clock), .in1(R6260));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6521 (.out1(R6522), .clock(clock), .in1(R6521));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6726 (.out1(R6727), .clock(clock), .in1(R6726));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6926 (.out1(R6927), .clock(clock), .in1(R6926));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7173 (.out1(R7174), .clock(clock), .in1(R7173));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7365 (.out1(R7366), .clock(clock), .in1(R7365));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7552 (.out1(R7553), .clock(clock), .in1(R7552));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7786 (.out1(R7787), .clock(clock), .in1(R7786));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7965 (.out1(R7966), .clock(clock), .in1(R7965));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8139 (.out1(R8140), .clock(clock), .in1(R8139));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8360 (.out1(R8361), .clock(clock), .in1(R8360));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8526 (.out1(R8527), .clock(clock), .in1(R8526));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8687 (.out1(R8688), .clock(clock), .in1(R8687));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8895 (.out1(R8896), .clock(clock), .in1(R8895));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9048 (.out1(R9049), .clock(clock), .in1(R9048));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9196 (.out1(R9197), .clock(clock), .in1(R9196));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9391 (.out1(R9392), .clock(clock), .in1(R9391));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9531 (.out1(R9532), .clock(clock), .in1(R9531));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9666 (.out1(R9667), .clock(clock), .in1(R9666));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9848 (.out1(R9849), .clock(clock), .in1(R9848));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9975 (.out1(R9976), .clock(clock), .in1(R9975));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10097 (.out1(R10098), .clock(clock), .in1(R10097));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10229 (.out1(R10230), .clock(clock), .in1(_944));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10230 (.out1(R10231), .clock(clock), .in1(_916));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10231 (.out1(R10232), .clock(clock), .in1(_896));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10232 (.out1(R10233), .clock(clock), .in1(_885));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10233 (.out1(R10234), .clock(clock), .in1(_878));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10234 (.out1(R10235), .clock(clock), .in1(_942));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10235 (.out1(R10236), .clock(clock), .in1(_935));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10236 (.out1(R10237), .clock(clock), .in1(_924));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10237 (.out1(R10238), .clock(clock), .in1(_904));
  SRAM op974 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_943),.ADR(R10235));
  SRAM op967 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_936),.ADR(R10236));
  SRAM op956 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_925),.ADR(R10237));
  SRAM op936 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_905),.ADR(R10238));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op968 (.out1(_937), .in1(2 'd 2), .in2(R9976));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op957 (.out1(_926), .in1(2 'd 2), .in2(R9976));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op950 (.out1(_919), .in1(2 'd 2), .in2(R9976));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op937 (.out1(_906), .in1(2 'd 2), .in2(R9976));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op930 (.out1(_899), .in1(2 'd 2), .in2(R9976));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op919 (.out1(_888), .in1(2 'd 2), .in2(R9976));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op948 (.out1(_917), .in1(vec70_3612_D), .in2(R10231));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op928 (.out1(_897), .in1(vec70_3612_D), .in2(R10232));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op917 (.out1(_886), .in1(vec70_3612_D), .in2(R10233));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op910 (.out1(_879), .in1(vec70_3612_D), .in2(R10234));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op976 (.out1(_945), .in1(R10230), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3814 (.out1(R3815), .clock(clock), .in1(R3814));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4070 (.out1(R4071), .clock(clock), .in1(R4070));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4325 (.out1(R4326), .clock(clock), .in1(R4325));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4570 (.out1(R4571), .clock(clock), .in1(R4570));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4810 (.out1(R4811), .clock(clock), .in1(R4810));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5097 (.out1(R5098), .clock(clock), .in1(R5097));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5329 (.out1(R5330), .clock(clock), .in1(R5329));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5556 (.out1(R5557), .clock(clock), .in1(R5556));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5830 (.out1(R5831), .clock(clock), .in1(R5830));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6048 (.out1(R6049), .clock(clock), .in1(R6048));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6261 (.out1(R6262), .clock(clock), .in1(R6261));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6522 (.out1(R6523), .clock(clock), .in1(R6522));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6727 (.out1(R6728), .clock(clock), .in1(R6727));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6927 (.out1(R6928), .clock(clock), .in1(R6927));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7174 (.out1(R7175), .clock(clock), .in1(R7174));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7366 (.out1(R7367), .clock(clock), .in1(R7366));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7553 (.out1(R7554), .clock(clock), .in1(R7553));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7787 (.out1(R7788), .clock(clock), .in1(R7787));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7966 (.out1(R7967), .clock(clock), .in1(R7966));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8140 (.out1(R8141), .clock(clock), .in1(R8140));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8361 (.out1(R8362), .clock(clock), .in1(R8361));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8527 (.out1(R8528), .clock(clock), .in1(R8527));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8688 (.out1(R8689), .clock(clock), .in1(R8688));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8896 (.out1(R8897), .clock(clock), .in1(R8896));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9049 (.out1(R9050), .clock(clock), .in1(R9049));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9197 (.out1(R9198), .clock(clock), .in1(R9197));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9392 (.out1(R9393), .clock(clock), .in1(R9392));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9532 (.out1(R9533), .clock(clock), .in1(R9532));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9667 (.out1(R9668), .clock(clock), .in1(R9667));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9849 (.out1(R9850), .clock(clock), .in1(R9849));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9976 (.out1(R9977), .clock(clock), .in1(R9976));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10098 (.out1(R10099), .clock(clock), .in1(R10098));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10238 (.out1(R10239), .clock(clock), .in1(_943));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10239 (.out1(R10240), .clock(clock), .in1(_936));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10240 (.out1(R10241), .clock(clock), .in1(_925));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10241 (.out1(R10242), .clock(clock), .in1(_905));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10242 (.out1(R10243), .clock(clock), .in1(_937));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10243 (.out1(R10244), .clock(clock), .in1(_926));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10244 (.out1(R10245), .clock(clock), .in1(_919));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10245 (.out1(R10246), .clock(clock), .in1(_906));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10246 (.out1(R10247), .clock(clock), .in1(_899));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10247 (.out1(R10248), .clock(clock), .in1(_888));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10248 (.out1(R10249), .clock(clock), .in1(_917));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10249 (.out1(R10250), .clock(clock), .in1(_897));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10250 (.out1(R10251), .clock(clock), .in1(_886));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10251 (.out1(R10252), .clock(clock), .in1(_879));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10252 (.out1(R10253), .clock(clock), .in1(_945));
  SRAM op949 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_918),.ADR(R10249));
  SRAM op929 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_898),.ADR(R10250));
  SRAM op918 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_887),.ADR(R10251));
  SRAM op911 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_880),.ADR(R10252));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op977 (.out1(_946), .in1(R10239), .in2(R10253));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op978 (.out1(_947), .in1(_946), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op969 (.out1(_938), .in1(R10243), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op958 (.out1(_927), .in1(R10244), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op938 (.out1(_907), .in1(R10246), .in2(64 'd 18446744073709551615));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op912 (.out1(_881), .in1(2 'd 2), .in2(R9977));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op979 (.out1(_948), .in1(_947), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op970 (.out1(_939), .in1(R10240), .in2(_938));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op959 (.out1(_928), .in1(R10241), .in2(_927));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op939 (.out1(_908), .in1(R10242), .in2(_907));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op980 (.out1(_949), .in1(_939), .in2(_948));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op960 (.out1(_929), .in1(_928), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op951 (.out1(_920), .in1(R10245), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op940 (.out1(_909), .in1(_908), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op931 (.out1(_900), .in1(R10247), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op920 (.out1(_889), .in1(R10248), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3815 (.out1(R3816), .clock(clock), .in1(R3815));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4071 (.out1(R4072), .clock(clock), .in1(R4071));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4326 (.out1(R4327), .clock(clock), .in1(R4326));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4571 (.out1(R4572), .clock(clock), .in1(R4571));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4811 (.out1(R4812), .clock(clock), .in1(R4811));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5098 (.out1(R5099), .clock(clock), .in1(R5098));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5330 (.out1(R5331), .clock(clock), .in1(R5330));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5557 (.out1(R5558), .clock(clock), .in1(R5557));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5831 (.out1(R5832), .clock(clock), .in1(R5831));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6049 (.out1(R6050), .clock(clock), .in1(R6049));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6262 (.out1(R6263), .clock(clock), .in1(R6262));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6523 (.out1(R6524), .clock(clock), .in1(R6523));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6728 (.out1(R6729), .clock(clock), .in1(R6728));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6928 (.out1(R6929), .clock(clock), .in1(R6928));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7175 (.out1(R7176), .clock(clock), .in1(R7175));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7367 (.out1(R7368), .clock(clock), .in1(R7367));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7554 (.out1(R7555), .clock(clock), .in1(R7554));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7788 (.out1(R7789), .clock(clock), .in1(R7788));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7967 (.out1(R7968), .clock(clock), .in1(R7967));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8141 (.out1(R8142), .clock(clock), .in1(R8141));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8362 (.out1(R8363), .clock(clock), .in1(R8362));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8528 (.out1(R8529), .clock(clock), .in1(R8528));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8689 (.out1(R8690), .clock(clock), .in1(R8689));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8897 (.out1(R8898), .clock(clock), .in1(R8897));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9050 (.out1(R9051), .clock(clock), .in1(R9050));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9198 (.out1(R9199), .clock(clock), .in1(R9198));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9393 (.out1(R9394), .clock(clock), .in1(R9393));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9533 (.out1(R9534), .clock(clock), .in1(R9533));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9668 (.out1(R9669), .clock(clock), .in1(R9668));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9850 (.out1(R9851), .clock(clock), .in1(R9850));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9977 (.out1(R9978), .clock(clock), .in1(R9977));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10099 (.out1(R10100), .clock(clock), .in1(R10099));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10253 (.out1(R10254), .clock(clock), .in1(_918));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10254 (.out1(R10255), .clock(clock), .in1(_898));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10255 (.out1(R10256), .clock(clock), .in1(_887));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10256 (.out1(R10257), .clock(clock), .in1(_880));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10257 (.out1(R10258), .clock(clock), .in1(_881));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10258 (.out1(R10259), .clock(clock), .in1(_949));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10259 (.out1(R10260), .clock(clock), .in1(_929));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10260 (.out1(R10261), .clock(clock), .in1(_920));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10261 (.out1(R10262), .clock(clock), .in1(_909));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10262 (.out1(R10263), .clock(clock), .in1(_900));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10263 (.out1(R10264), .clock(clock), .in1(_889));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op961 (.out1(_930), .in1(R10260), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op952 (.out1(_921), .in1(R10254), .in2(R10261));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op921 (.out1(_890), .in1(R10256), .in2(R10264));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op981 (.out1(_950), .in1(R10259), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op962 (.out1(_931), .in1(_921), .in2(_930));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op941 (.out1(_910), .in1(R10262), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op932 (.out1(_901), .in1(R10255), .in2(R10263));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op922 (.out1(_891), .in1(_890), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op913 (.out1(_882), .in1(R10258), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op942 (.out1(_911), .in1(_901), .in2(_910));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op982 (.out1(_951), .in1(_950), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op963 (.out1(_932), .in1(_931), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op923 (.out1(_892), .in1(_891), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op914 (.out1(_883), .in1(R10257), .in2(_882));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op983 (.out1(_952), .in1(_932), .in2(_951));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op943 (.out1(_912), .in1(_911), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op924 (.out1(_893), .in1(_883), .in2(_892));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3816 (.out1(R3817), .clock(clock), .in1(R3816));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4072 (.out1(R4073), .clock(clock), .in1(R4072));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4327 (.out1(R4328), .clock(clock), .in1(R4327));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4572 (.out1(R4573), .clock(clock), .in1(R4572));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4812 (.out1(R4813), .clock(clock), .in1(R4812));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5099 (.out1(R5100), .clock(clock), .in1(R5099));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5331 (.out1(R5332), .clock(clock), .in1(R5331));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5558 (.out1(R5559), .clock(clock), .in1(R5558));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5832 (.out1(R5833), .clock(clock), .in1(R5832));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6050 (.out1(R6051), .clock(clock), .in1(R6050));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6263 (.out1(R6264), .clock(clock), .in1(R6263));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6524 (.out1(R6525), .clock(clock), .in1(R6524));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6729 (.out1(R6730), .clock(clock), .in1(R6729));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6929 (.out1(R6930), .clock(clock), .in1(R6929));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7176 (.out1(R7177), .clock(clock), .in1(R7176));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7368 (.out1(R7369), .clock(clock), .in1(R7368));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7555 (.out1(R7556), .clock(clock), .in1(R7555));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7789 (.out1(R7790), .clock(clock), .in1(R7789));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7968 (.out1(R7969), .clock(clock), .in1(R7968));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8142 (.out1(R8143), .clock(clock), .in1(R8142));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8363 (.out1(R8364), .clock(clock), .in1(R8363));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8529 (.out1(R8530), .clock(clock), .in1(R8529));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8690 (.out1(R8691), .clock(clock), .in1(R8690));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8898 (.out1(R8899), .clock(clock), .in1(R8898));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9051 (.out1(R9052), .clock(clock), .in1(R9051));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9199 (.out1(R9200), .clock(clock), .in1(R9199));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9394 (.out1(R9395), .clock(clock), .in1(R9394));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9534 (.out1(R9535), .clock(clock), .in1(R9534));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9669 (.out1(R9670), .clock(clock), .in1(R9669));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9851 (.out1(R9852), .clock(clock), .in1(R9851));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9978 (.out1(R9979), .clock(clock), .in1(R9978));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10100 (.out1(R10101), .clock(clock), .in1(R10100));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10264 (.out1(R10265), .clock(clock), .in1(_952));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10265 (.out1(R10266), .clock(clock), .in1(_912));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10266 (.out1(R10267), .clock(clock), .in1(_893));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op904 (.out1(_873), .in1(R9852));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op944 (.out1(_913), .in1(R10266), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op925 (.out1(_894), .in1(R10267), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op984 (.out1(_953), .in1(R10265), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op945 (.out1(_914), .in1(_894), .in2(_913));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op905 (.out1(_874), .in1(_873), .in2(2 'd 2));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op985 (.out1(_954), .in1(_914), .in2(_953));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op986 (.out1(_955), .in1(_954), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3817 (.out1(R3818), .clock(clock), .in1(R3817));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4073 (.out1(R4074), .clock(clock), .in1(R4073));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4328 (.out1(R4329), .clock(clock), .in1(R4328));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4573 (.out1(R4574), .clock(clock), .in1(R4573));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4813 (.out1(R4814), .clock(clock), .in1(R4813));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5100 (.out1(R5101), .clock(clock), .in1(R5100));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5332 (.out1(R5333), .clock(clock), .in1(R5332));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5559 (.out1(R5560), .clock(clock), .in1(R5559));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5833 (.out1(R5834), .clock(clock), .in1(R5833));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6051 (.out1(R6052), .clock(clock), .in1(R6051));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6264 (.out1(R6265), .clock(clock), .in1(R6264));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6525 (.out1(R6526), .clock(clock), .in1(R6525));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6730 (.out1(R6731), .clock(clock), .in1(R6730));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6930 (.out1(R6931), .clock(clock), .in1(R6930));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7177 (.out1(R7178), .clock(clock), .in1(R7177));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7369 (.out1(R7370), .clock(clock), .in1(R7369));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7556 (.out1(R7557), .clock(clock), .in1(R7556));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7790 (.out1(R7791), .clock(clock), .in1(R7790));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7969 (.out1(R7970), .clock(clock), .in1(R7969));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8143 (.out1(R8144), .clock(clock), .in1(R8143));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8364 (.out1(R8365), .clock(clock), .in1(R8364));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8530 (.out1(R8531), .clock(clock), .in1(R8530));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8691 (.out1(R8692), .clock(clock), .in1(R8691));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8899 (.out1(R8900), .clock(clock), .in1(R8899));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9052 (.out1(R9053), .clock(clock), .in1(R9052));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9200 (.out1(R9201), .clock(clock), .in1(R9200));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9395 (.out1(R9396), .clock(clock), .in1(R9395));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9535 (.out1(R9536), .clock(clock), .in1(R9535));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9670 (.out1(R9671), .clock(clock), .in1(R9670));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9852 (.out1(R9853), .clock(clock), .in1(R9852));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9979 (.out1(R9980), .clock(clock), .in1(R9979));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10101 (.out1(R10102), .clock(clock), .in1(R10101));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10267 (.out1(R10268), .clock(clock), .in1(_874));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10268 (.out1(R10269), .clock(clock), .in1(_955));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op987 (.out1(_956), .in1(R10269), .in2(57 'd 72340172838076673));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op906 (.out1(_875), .in1(base0_70_3617_D), .in2(R10268));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3818 (.out1(R3819), .clock(clock), .in1(R3818));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4074 (.out1(R4075), .clock(clock), .in1(R4074));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4329 (.out1(R4330), .clock(clock), .in1(R4329));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4574 (.out1(R4575), .clock(clock), .in1(R4574));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4814 (.out1(R4815), .clock(clock), .in1(R4814));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5101 (.out1(R5102), .clock(clock), .in1(R5101));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5333 (.out1(R5334), .clock(clock), .in1(R5333));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5560 (.out1(R5561), .clock(clock), .in1(R5560));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5834 (.out1(R5835), .clock(clock), .in1(R5834));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6052 (.out1(R6053), .clock(clock), .in1(R6052));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6265 (.out1(R6266), .clock(clock), .in1(R6265));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6526 (.out1(R6527), .clock(clock), .in1(R6526));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6731 (.out1(R6732), .clock(clock), .in1(R6731));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6931 (.out1(R6932), .clock(clock), .in1(R6931));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7178 (.out1(R7179), .clock(clock), .in1(R7178));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7370 (.out1(R7371), .clock(clock), .in1(R7370));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7557 (.out1(R7558), .clock(clock), .in1(R7557));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7791 (.out1(R7792), .clock(clock), .in1(R7791));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7970 (.out1(R7971), .clock(clock), .in1(R7970));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8144 (.out1(R8145), .clock(clock), .in1(R8144));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8365 (.out1(R8366), .clock(clock), .in1(R8365));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8531 (.out1(R8532), .clock(clock), .in1(R8531));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8692 (.out1(R8693), .clock(clock), .in1(R8692));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8900 (.out1(R8901), .clock(clock), .in1(R8900));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9053 (.out1(R9054), .clock(clock), .in1(R9053));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9201 (.out1(R9202), .clock(clock), .in1(R9201));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9396 (.out1(R9397), .clock(clock), .in1(R9396));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9536 (.out1(R9537), .clock(clock), .in1(R9536));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9671 (.out1(R9672), .clock(clock), .in1(R9671));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9853 (.out1(R9854), .clock(clock), .in1(R9853));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9980 (.out1(R9981), .clock(clock), .in1(R9980));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10102 (.out1(R10103), .clock(clock), .in1(R10102));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10269 (.out1(R10270), .clock(clock), .in1(_956));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10270 (.out1(R10271), .clock(clock), .in1(_875));
  SRAM op907 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_876),.ADR(R10271));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op988 (.out1(_957), .in1(R10270), .in2(6 'd 56));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3819 (.out1(R3820), .clock(clock), .in1(R3819));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4075 (.out1(R4076), .clock(clock), .in1(R4075));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4330 (.out1(R4331), .clock(clock), .in1(R4330));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4575 (.out1(R4576), .clock(clock), .in1(R4575));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4815 (.out1(R4816), .clock(clock), .in1(R4815));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5102 (.out1(R5103), .clock(clock), .in1(R5102));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5334 (.out1(R5335), .clock(clock), .in1(R5334));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5561 (.out1(R5562), .clock(clock), .in1(R5561));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5835 (.out1(R5836), .clock(clock), .in1(R5835));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6053 (.out1(R6054), .clock(clock), .in1(R6053));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6266 (.out1(R6267), .clock(clock), .in1(R6266));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6527 (.out1(R6528), .clock(clock), .in1(R6527));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6732 (.out1(R6733), .clock(clock), .in1(R6732));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6932 (.out1(R6933), .clock(clock), .in1(R6932));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7179 (.out1(R7180), .clock(clock), .in1(R7179));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7371 (.out1(R7372), .clock(clock), .in1(R7371));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7558 (.out1(R7559), .clock(clock), .in1(R7558));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7792 (.out1(R7793), .clock(clock), .in1(R7792));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7971 (.out1(R7972), .clock(clock), .in1(R7971));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8145 (.out1(R8146), .clock(clock), .in1(R8145));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8366 (.out1(R8367), .clock(clock), .in1(R8366));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8532 (.out1(R8533), .clock(clock), .in1(R8532));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8693 (.out1(R8694), .clock(clock), .in1(R8693));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8901 (.out1(R8902), .clock(clock), .in1(R8901));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9054 (.out1(R9055), .clock(clock), .in1(R9054));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9202 (.out1(R9203), .clock(clock), .in1(R9202));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9397 (.out1(R9398), .clock(clock), .in1(R9397));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9537 (.out1(R9538), .clock(clock), .in1(R9537));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9672 (.out1(R9673), .clock(clock), .in1(R9672));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9854 (.out1(R9855), .clock(clock), .in1(R9854));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9981 (.out1(R9982), .clock(clock), .in1(R9981));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10103 (.out1(R10104), .clock(clock), .in1(R10103));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10271 (.out1(R10272), .clock(clock), .in1(_876));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10272 (.out1(R10273), .clock(clock), .in1(_957));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op989 (.out1(_958), .in1(R10273));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op990 (.out1(_959), .in1(R10272), .in2(_958));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op991 (.out1(idx_3618), .in1(_959), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3820 (.out1(R3821), .clock(clock), .in1(R3820));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4076 (.out1(R4077), .clock(clock), .in1(R4076));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4331 (.out1(R4332), .clock(clock), .in1(R4331));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4576 (.out1(R4577), .clock(clock), .in1(R4576));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4816 (.out1(R4817), .clock(clock), .in1(R4816));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5103 (.out1(R5104), .clock(clock), .in1(R5103));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5335 (.out1(R5336), .clock(clock), .in1(R5335));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5562 (.out1(R5563), .clock(clock), .in1(R5562));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5836 (.out1(R5837), .clock(clock), .in1(R5836));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6054 (.out1(R6055), .clock(clock), .in1(R6054));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6267 (.out1(R6268), .clock(clock), .in1(R6267));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6528 (.out1(R6529), .clock(clock), .in1(R6528));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6733 (.out1(R6734), .clock(clock), .in1(R6733));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6933 (.out1(R6934), .clock(clock), .in1(R6933));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7180 (.out1(R7181), .clock(clock), .in1(R7180));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7372 (.out1(R7373), .clock(clock), .in1(R7372));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7559 (.out1(R7560), .clock(clock), .in1(R7559));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7793 (.out1(R7794), .clock(clock), .in1(R7793));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7972 (.out1(R7973), .clock(clock), .in1(R7972));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8146 (.out1(R8147), .clock(clock), .in1(R8146));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8367 (.out1(R8368), .clock(clock), .in1(R8367));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8533 (.out1(R8534), .clock(clock), .in1(R8533));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8694 (.out1(R8695), .clock(clock), .in1(R8694));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8902 (.out1(R8903), .clock(clock), .in1(R8902));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9055 (.out1(R9056), .clock(clock), .in1(R9055));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9203 (.out1(R9204), .clock(clock), .in1(R9203));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9398 (.out1(R9399), .clock(clock), .in1(R9398));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9538 (.out1(R9539), .clock(clock), .in1(R9538));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9673 (.out1(R9674), .clock(clock), .in1(R9673));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9855 (.out1(R9856), .clock(clock), .in1(R9855));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9982 (.out1(R9983), .clock(clock), .in1(R9982));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10104 (.out1(R10105), .clock(clock), .in1(R10104));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10273 (.out1(R10274), .clock(clock), .in1(idx_3618));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op995 (.out1(_962), .in1(R10274));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op996 (.out1(_963), .in1(_962), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3821 (.out1(R3822), .clock(clock), .in1(R3821));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4077 (.out1(R4078), .clock(clock), .in1(R4077));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4332 (.out1(R4333), .clock(clock), .in1(R4332));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4577 (.out1(R4578), .clock(clock), .in1(R4577));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4817 (.out1(R4818), .clock(clock), .in1(R4817));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5104 (.out1(R5105), .clock(clock), .in1(R5104));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5336 (.out1(R5337), .clock(clock), .in1(R5336));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5563 (.out1(R5564), .clock(clock), .in1(R5563));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5837 (.out1(R5838), .clock(clock), .in1(R5837));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6055 (.out1(R6056), .clock(clock), .in1(R6055));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6268 (.out1(R6269), .clock(clock), .in1(R6268));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6529 (.out1(R6530), .clock(clock), .in1(R6529));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6734 (.out1(R6735), .clock(clock), .in1(R6734));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6934 (.out1(R6935), .clock(clock), .in1(R6934));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7181 (.out1(R7182), .clock(clock), .in1(R7181));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7373 (.out1(R7374), .clock(clock), .in1(R7373));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7560 (.out1(R7561), .clock(clock), .in1(R7560));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7794 (.out1(R7795), .clock(clock), .in1(R7794));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7973 (.out1(R7974), .clock(clock), .in1(R7973));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8147 (.out1(R8148), .clock(clock), .in1(R8147));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8368 (.out1(R8369), .clock(clock), .in1(R8368));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8534 (.out1(R8535), .clock(clock), .in1(R8534));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8695 (.out1(R8696), .clock(clock), .in1(R8695));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8903 (.out1(R8904), .clock(clock), .in1(R8903));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9056 (.out1(R9057), .clock(clock), .in1(R9056));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9204 (.out1(R9205), .clock(clock), .in1(R9204));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9399 (.out1(R9400), .clock(clock), .in1(R9399));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9539 (.out1(R9540), .clock(clock), .in1(R9539));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9674 (.out1(R9675), .clock(clock), .in1(R9674));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9856 (.out1(R9857), .clock(clock), .in1(R9856));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9983 (.out1(R9984), .clock(clock), .in1(R9983));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10105 (.out1(R10106), .clock(clock), .in1(R10105));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10274 (.out1(R10275), .clock(clock), .in1(R10274));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10387 (.out1(R10388), .clock(clock), .in1(_963));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op997 (.out1(_964), .in1(vec76_3620_D), .in2(R10388));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3822 (.out1(R3823), .clock(clock), .in1(R3822));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4078 (.out1(R4079), .clock(clock), .in1(R4078));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4333 (.out1(R4334), .clock(clock), .in1(R4333));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4578 (.out1(R4579), .clock(clock), .in1(R4578));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4818 (.out1(R4819), .clock(clock), .in1(R4818));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5105 (.out1(R5106), .clock(clock), .in1(R5105));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5337 (.out1(R5338), .clock(clock), .in1(R5337));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5564 (.out1(R5565), .clock(clock), .in1(R5564));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5838 (.out1(R5839), .clock(clock), .in1(R5838));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6056 (.out1(R6057), .clock(clock), .in1(R6056));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6269 (.out1(R6270), .clock(clock), .in1(R6269));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6530 (.out1(R6531), .clock(clock), .in1(R6530));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6735 (.out1(R6736), .clock(clock), .in1(R6735));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6935 (.out1(R6936), .clock(clock), .in1(R6935));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7182 (.out1(R7183), .clock(clock), .in1(R7182));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7374 (.out1(R7375), .clock(clock), .in1(R7374));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7561 (.out1(R7562), .clock(clock), .in1(R7561));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7795 (.out1(R7796), .clock(clock), .in1(R7795));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7974 (.out1(R7975), .clock(clock), .in1(R7974));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8148 (.out1(R8149), .clock(clock), .in1(R8148));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8369 (.out1(R8370), .clock(clock), .in1(R8369));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8535 (.out1(R8536), .clock(clock), .in1(R8535));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8696 (.out1(R8697), .clock(clock), .in1(R8696));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8904 (.out1(R8905), .clock(clock), .in1(R8904));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9057 (.out1(R9058), .clock(clock), .in1(R9057));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9205 (.out1(R9206), .clock(clock), .in1(R9205));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9400 (.out1(R9401), .clock(clock), .in1(R9400));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9540 (.out1(R9541), .clock(clock), .in1(R9540));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9675 (.out1(R9676), .clock(clock), .in1(R9675));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9857 (.out1(R9858), .clock(clock), .in1(R9857));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9984 (.out1(R9985), .clock(clock), .in1(R9984));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10106 (.out1(R10107), .clock(clock), .in1(R10106));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10275 (.out1(R10276), .clock(clock), .in1(R10275));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10388 (.out1(R10389), .clock(clock), .in1(_964));
  SRAM op998 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_965),.ADR(R10389));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3823 (.out1(R3824), .clock(clock), .in1(R3823));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4079 (.out1(R4080), .clock(clock), .in1(R4079));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4334 (.out1(R4335), .clock(clock), .in1(R4334));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4579 (.out1(R4580), .clock(clock), .in1(R4579));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4819 (.out1(R4820), .clock(clock), .in1(R4819));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5106 (.out1(R5107), .clock(clock), .in1(R5106));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5338 (.out1(R5339), .clock(clock), .in1(R5338));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5565 (.out1(R5566), .clock(clock), .in1(R5565));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5839 (.out1(R5840), .clock(clock), .in1(R5839));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6057 (.out1(R6058), .clock(clock), .in1(R6057));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6270 (.out1(R6271), .clock(clock), .in1(R6270));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6531 (.out1(R6532), .clock(clock), .in1(R6531));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6736 (.out1(R6737), .clock(clock), .in1(R6736));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6936 (.out1(R6937), .clock(clock), .in1(R6936));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7183 (.out1(R7184), .clock(clock), .in1(R7183));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7375 (.out1(R7376), .clock(clock), .in1(R7375));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7562 (.out1(R7563), .clock(clock), .in1(R7562));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7796 (.out1(R7797), .clock(clock), .in1(R7796));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7975 (.out1(R7976), .clock(clock), .in1(R7975));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8149 (.out1(R8150), .clock(clock), .in1(R8149));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8370 (.out1(R8371), .clock(clock), .in1(R8370));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8536 (.out1(R8537), .clock(clock), .in1(R8536));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8697 (.out1(R8698), .clock(clock), .in1(R8697));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8905 (.out1(R8906), .clock(clock), .in1(R8905));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9058 (.out1(R9059), .clock(clock), .in1(R9058));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9206 (.out1(R9207), .clock(clock), .in1(R9206));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9401 (.out1(R9402), .clock(clock), .in1(R9401));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9541 (.out1(R9542), .clock(clock), .in1(R9541));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9676 (.out1(R9677), .clock(clock), .in1(R9676));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9858 (.out1(R9859), .clock(clock), .in1(R9858));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9985 (.out1(R9986), .clock(clock), .in1(R9985));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10107 (.out1(R10108), .clock(clock), .in1(R10107));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10276 (.out1(R10277), .clock(clock), .in1(R10276));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10389 (.out1(R10390), .clock(clock), .in1(_965));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op992 (.out1(_960), .in1(ip2_3602_D), .in2(6 'd 46));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op993 (.out1(_961), .in1(_960));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op994 (.out1(off_3619), .in1(_961), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op999 (.out1(_966), .in1(R10390), .in2(off_3619));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3824 (.out1(R3825), .clock(clock), .in1(R3824));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4080 (.out1(R4081), .clock(clock), .in1(R4080));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4335 (.out1(R4336), .clock(clock), .in1(R4335));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4580 (.out1(R4581), .clock(clock), .in1(R4580));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4820 (.out1(R4821), .clock(clock), .in1(R4820));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5107 (.out1(R5108), .clock(clock), .in1(R5107));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5339 (.out1(R5340), .clock(clock), .in1(R5339));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5566 (.out1(R5567), .clock(clock), .in1(R5566));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5840 (.out1(R5841), .clock(clock), .in1(R5840));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6058 (.out1(R6059), .clock(clock), .in1(R6058));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6271 (.out1(R6272), .clock(clock), .in1(R6271));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6532 (.out1(R6533), .clock(clock), .in1(R6532));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6737 (.out1(R6738), .clock(clock), .in1(R6737));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6937 (.out1(R6938), .clock(clock), .in1(R6937));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7184 (.out1(R7185), .clock(clock), .in1(R7184));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7376 (.out1(R7377), .clock(clock), .in1(R7376));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7563 (.out1(R7564), .clock(clock), .in1(R7563));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7797 (.out1(R7798), .clock(clock), .in1(R7797));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7976 (.out1(R7977), .clock(clock), .in1(R7976));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8150 (.out1(R8151), .clock(clock), .in1(R8150));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8371 (.out1(R8372), .clock(clock), .in1(R8371));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8537 (.out1(R8538), .clock(clock), .in1(R8537));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8698 (.out1(R8699), .clock(clock), .in1(R8698));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8906 (.out1(R8907), .clock(clock), .in1(R8906));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9059 (.out1(R9060), .clock(clock), .in1(R9059));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9207 (.out1(R9208), .clock(clock), .in1(R9207));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9402 (.out1(R9403), .clock(clock), .in1(R9402));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9542 (.out1(R9543), .clock(clock), .in1(R9542));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9677 (.out1(R9678), .clock(clock), .in1(R9677));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9859 (.out1(R9860), .clock(clock), .in1(R9859));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9986 (.out1(R9987), .clock(clock), .in1(R9986));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10108 (.out1(R10109), .clock(clock), .in1(R10108));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10277 (.out1(R10278), .clock(clock), .in1(R10277));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10390 (.out1(R10391), .clock(clock), .in1(off_3619));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10498 (.out1(R10499), .clock(clock), .in1(_966));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op1000 (.out1(_967), .in1(R10499), .in2(1 'd 1));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op1001 (.out1(ifout1001), .in1(_967), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1069 (.out1(_1035), .in1(R10278));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1062 (.out1(_1028), .in1(R10278));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1051 (.out1(_1017), .in1(R10278));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1031 (.out1(_997), .in1(R10278));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1070 (.out1(_1036), .in1(_1035), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1063 (.out1(_1029), .in1(_1028), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1052 (.out1(_1018), .in1(_1017), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1032 (.out1(_998), .in1(_997), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3825 (.out1(R3826), .clock(clock), .in1(R3825));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4081 (.out1(R4082), .clock(clock), .in1(R4081));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4336 (.out1(R4337), .clock(clock), .in1(R4336));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4581 (.out1(R4582), .clock(clock), .in1(R4581));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4821 (.out1(R4822), .clock(clock), .in1(R4821));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5108 (.out1(R5109), .clock(clock), .in1(R5108));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5340 (.out1(R5341), .clock(clock), .in1(R5340));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5567 (.out1(R5568), .clock(clock), .in1(R5567));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5841 (.out1(R5842), .clock(clock), .in1(R5841));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6059 (.out1(R6060), .clock(clock), .in1(R6059));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6272 (.out1(R6273), .clock(clock), .in1(R6272));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6533 (.out1(R6534), .clock(clock), .in1(R6533));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6738 (.out1(R6739), .clock(clock), .in1(R6738));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6938 (.out1(R6939), .clock(clock), .in1(R6938));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7185 (.out1(R7186), .clock(clock), .in1(R7185));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7377 (.out1(R7378), .clock(clock), .in1(R7377));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7564 (.out1(R7565), .clock(clock), .in1(R7564));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7798 (.out1(R7799), .clock(clock), .in1(R7798));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7977 (.out1(R7978), .clock(clock), .in1(R7977));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8151 (.out1(R8152), .clock(clock), .in1(R8151));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8372 (.out1(R8373), .clock(clock), .in1(R8372));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8538 (.out1(R8539), .clock(clock), .in1(R8538));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8699 (.out1(R8700), .clock(clock), .in1(R8699));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8907 (.out1(R8908), .clock(clock), .in1(R8907));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9060 (.out1(R9061), .clock(clock), .in1(R9060));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9208 (.out1(R9209), .clock(clock), .in1(R9208));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9403 (.out1(R9404), .clock(clock), .in1(R9403));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9543 (.out1(R9544), .clock(clock), .in1(R9543));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9678 (.out1(R9679), .clock(clock), .in1(R9678));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9860 (.out1(R9861), .clock(clock), .in1(R9860));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9987 (.out1(R9988), .clock(clock), .in1(R9987));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10109 (.out1(R10110), .clock(clock), .in1(R10109));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10278 (.out1(R10279), .clock(clock), .in1(R10278));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10391 (.out1(R10392), .clock(clock), .in1(R10391));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10499 (.out1(R10500), .clock(clock), .in1(ifout1001));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10615 (.out1(R10616), .clock(clock), .in1(_1036));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10616 (.out1(R10617), .clock(clock), .in1(_1029));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10617 (.out1(R10618), .clock(clock), .in1(_1018));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10618 (.out1(R10619), .clock(clock), .in1(_998));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1044 (.out1(_1010), .in1(R10279));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1024 (.out1(_990), .in1(R10279));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1013 (.out1(_979), .in1(R10279));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1006 (.out1(_972), .in1(R10279));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1073 (.out1(_1039), .in1(2 'd 2), .in2(R10392));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1045 (.out1(_1011), .in1(_1010), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1025 (.out1(_991), .in1(_990), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1014 (.out1(_980), .in1(_979), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1007 (.out1(_973), .in1(_972), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1071 (.out1(_1037), .in1(vec76_3620_D), .in2(R10616));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1064 (.out1(_1030), .in1(vec76_3620_D), .in2(R10617));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1053 (.out1(_1019), .in1(vec76_3620_D), .in2(R10618));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1033 (.out1(_999), .in1(vec76_3620_D), .in2(R10619));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3826 (.out1(R3827), .clock(clock), .in1(R3826));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4082 (.out1(R4083), .clock(clock), .in1(R4082));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4337 (.out1(R4338), .clock(clock), .in1(R4337));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4582 (.out1(R4583), .clock(clock), .in1(R4582));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4822 (.out1(R4823), .clock(clock), .in1(R4822));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5109 (.out1(R5110), .clock(clock), .in1(R5109));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5341 (.out1(R5342), .clock(clock), .in1(R5341));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5568 (.out1(R5569), .clock(clock), .in1(R5568));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5842 (.out1(R5843), .clock(clock), .in1(R5842));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6060 (.out1(R6061), .clock(clock), .in1(R6060));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6273 (.out1(R6274), .clock(clock), .in1(R6273));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6534 (.out1(R6535), .clock(clock), .in1(R6534));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6739 (.out1(R6740), .clock(clock), .in1(R6739));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6939 (.out1(R6940), .clock(clock), .in1(R6939));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7186 (.out1(R7187), .clock(clock), .in1(R7186));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7378 (.out1(R7379), .clock(clock), .in1(R7378));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7565 (.out1(R7566), .clock(clock), .in1(R7565));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7799 (.out1(R7800), .clock(clock), .in1(R7799));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7978 (.out1(R7979), .clock(clock), .in1(R7978));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8152 (.out1(R8153), .clock(clock), .in1(R8152));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8373 (.out1(R8374), .clock(clock), .in1(R8373));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8539 (.out1(R8540), .clock(clock), .in1(R8539));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8700 (.out1(R8701), .clock(clock), .in1(R8700));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8908 (.out1(R8909), .clock(clock), .in1(R8908));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9061 (.out1(R9062), .clock(clock), .in1(R9061));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9209 (.out1(R9210), .clock(clock), .in1(R9209));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9404 (.out1(R9405), .clock(clock), .in1(R9404));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9544 (.out1(R9545), .clock(clock), .in1(R9544));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9679 (.out1(R9680), .clock(clock), .in1(R9679));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9861 (.out1(R9862), .clock(clock), .in1(R9861));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9988 (.out1(R9989), .clock(clock), .in1(R9988));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10110 (.out1(R10111), .clock(clock), .in1(R10110));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10279 (.out1(R10280), .clock(clock), .in1(R10279));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10392 (.out1(R10393), .clock(clock), .in1(R10392));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10500 (.out1(R10501), .clock(clock), .in1(R10500));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10619 (.out1(R10620), .clock(clock), .in1(_1039));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10620 (.out1(R10621), .clock(clock), .in1(_1011));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10621 (.out1(R10622), .clock(clock), .in1(_991));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10622 (.out1(R10623), .clock(clock), .in1(_980));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10623 (.out1(R10624), .clock(clock), .in1(_973));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10624 (.out1(R10625), .clock(clock), .in1(_1037));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10625 (.out1(R10626), .clock(clock), .in1(_1030));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10626 (.out1(R10627), .clock(clock), .in1(_1019));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10627 (.out1(R10628), .clock(clock), .in1(_999));
  SRAM op1072 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1038),.ADR(R10625));
  SRAM op1065 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1031),.ADR(R10626));
  SRAM op1054 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1020),.ADR(R10627));
  SRAM op1034 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1000),.ADR(R10628));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1066 (.out1(_1032), .in1(2 'd 2), .in2(R10393));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1055 (.out1(_1021), .in1(2 'd 2), .in2(R10393));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1048 (.out1(_1014), .in1(2 'd 2), .in2(R10393));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1035 (.out1(_1001), .in1(2 'd 2), .in2(R10393));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1028 (.out1(_994), .in1(2 'd 2), .in2(R10393));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1017 (.out1(_983), .in1(2 'd 2), .in2(R10393));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1046 (.out1(_1012), .in1(vec76_3620_D), .in2(R10621));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1026 (.out1(_992), .in1(vec76_3620_D), .in2(R10622));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1015 (.out1(_981), .in1(vec76_3620_D), .in2(R10623));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1008 (.out1(_974), .in1(vec76_3620_D), .in2(R10624));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1074 (.out1(_1040), .in1(R10620), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3827 (.out1(R3828), .clock(clock), .in1(R3827));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4083 (.out1(R4084), .clock(clock), .in1(R4083));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4338 (.out1(R4339), .clock(clock), .in1(R4338));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4583 (.out1(R4584), .clock(clock), .in1(R4583));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4823 (.out1(R4824), .clock(clock), .in1(R4823));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5110 (.out1(R5111), .clock(clock), .in1(R5110));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5342 (.out1(R5343), .clock(clock), .in1(R5342));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5569 (.out1(R5570), .clock(clock), .in1(R5569));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5843 (.out1(R5844), .clock(clock), .in1(R5843));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6061 (.out1(R6062), .clock(clock), .in1(R6061));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6274 (.out1(R6275), .clock(clock), .in1(R6274));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6535 (.out1(R6536), .clock(clock), .in1(R6535));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6740 (.out1(R6741), .clock(clock), .in1(R6740));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6940 (.out1(R6941), .clock(clock), .in1(R6940));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7187 (.out1(R7188), .clock(clock), .in1(R7187));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7379 (.out1(R7380), .clock(clock), .in1(R7379));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7566 (.out1(R7567), .clock(clock), .in1(R7566));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7800 (.out1(R7801), .clock(clock), .in1(R7800));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7979 (.out1(R7980), .clock(clock), .in1(R7979));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8153 (.out1(R8154), .clock(clock), .in1(R8153));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8374 (.out1(R8375), .clock(clock), .in1(R8374));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8540 (.out1(R8541), .clock(clock), .in1(R8540));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8701 (.out1(R8702), .clock(clock), .in1(R8701));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8909 (.out1(R8910), .clock(clock), .in1(R8909));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9062 (.out1(R9063), .clock(clock), .in1(R9062));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9210 (.out1(R9211), .clock(clock), .in1(R9210));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9405 (.out1(R9406), .clock(clock), .in1(R9405));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9545 (.out1(R9546), .clock(clock), .in1(R9545));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9680 (.out1(R9681), .clock(clock), .in1(R9680));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9862 (.out1(R9863), .clock(clock), .in1(R9862));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9989 (.out1(R9990), .clock(clock), .in1(R9989));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10111 (.out1(R10112), .clock(clock), .in1(R10111));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10280 (.out1(R10281), .clock(clock), .in1(R10280));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10393 (.out1(R10394), .clock(clock), .in1(R10393));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10501 (.out1(R10502), .clock(clock), .in1(R10501));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10628 (.out1(R10629), .clock(clock), .in1(_1038));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10629 (.out1(R10630), .clock(clock), .in1(_1031));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10630 (.out1(R10631), .clock(clock), .in1(_1020));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10631 (.out1(R10632), .clock(clock), .in1(_1000));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10632 (.out1(R10633), .clock(clock), .in1(_1032));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10633 (.out1(R10634), .clock(clock), .in1(_1021));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10634 (.out1(R10635), .clock(clock), .in1(_1014));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10635 (.out1(R10636), .clock(clock), .in1(_1001));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10636 (.out1(R10637), .clock(clock), .in1(_994));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10637 (.out1(R10638), .clock(clock), .in1(_983));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10638 (.out1(R10639), .clock(clock), .in1(_1012));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10639 (.out1(R10640), .clock(clock), .in1(_992));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10640 (.out1(R10641), .clock(clock), .in1(_981));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10641 (.out1(R10642), .clock(clock), .in1(_974));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10642 (.out1(R10643), .clock(clock), .in1(_1040));
  SRAM op1047 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1013),.ADR(R10639));
  SRAM op1027 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_993),.ADR(R10640));
  SRAM op1016 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_982),.ADR(R10641));
  SRAM op1009 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_975),.ADR(R10642));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1075 (.out1(_1041), .in1(R10629), .in2(R10643));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1076 (.out1(_1042), .in1(_1041), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1067 (.out1(_1033), .in1(R10633), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1056 (.out1(_1022), .in1(R10634), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1036 (.out1(_1002), .in1(R10636), .in2(64 'd 18446744073709551615));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1010 (.out1(_976), .in1(2 'd 2), .in2(R10394));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1077 (.out1(_1043), .in1(_1042), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1068 (.out1(_1034), .in1(R10630), .in2(_1033));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1057 (.out1(_1023), .in1(R10631), .in2(_1022));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1037 (.out1(_1003), .in1(R10632), .in2(_1002));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1078 (.out1(_1044), .in1(_1034), .in2(_1043));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1058 (.out1(_1024), .in1(_1023), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1049 (.out1(_1015), .in1(R10635), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1038 (.out1(_1004), .in1(_1003), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1029 (.out1(_995), .in1(R10637), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1018 (.out1(_984), .in1(R10638), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3828 (.out1(R3829), .clock(clock), .in1(R3828));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4084 (.out1(R4085), .clock(clock), .in1(R4084));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4339 (.out1(R4340), .clock(clock), .in1(R4339));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4584 (.out1(R4585), .clock(clock), .in1(R4584));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4824 (.out1(R4825), .clock(clock), .in1(R4824));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5111 (.out1(R5112), .clock(clock), .in1(R5111));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5343 (.out1(R5344), .clock(clock), .in1(R5343));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5570 (.out1(R5571), .clock(clock), .in1(R5570));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5844 (.out1(R5845), .clock(clock), .in1(R5844));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6062 (.out1(R6063), .clock(clock), .in1(R6062));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6275 (.out1(R6276), .clock(clock), .in1(R6275));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6536 (.out1(R6537), .clock(clock), .in1(R6536));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6741 (.out1(R6742), .clock(clock), .in1(R6741));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6941 (.out1(R6942), .clock(clock), .in1(R6941));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7188 (.out1(R7189), .clock(clock), .in1(R7188));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7380 (.out1(R7381), .clock(clock), .in1(R7380));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7567 (.out1(R7568), .clock(clock), .in1(R7567));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7801 (.out1(R7802), .clock(clock), .in1(R7801));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7980 (.out1(R7981), .clock(clock), .in1(R7980));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8154 (.out1(R8155), .clock(clock), .in1(R8154));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8375 (.out1(R8376), .clock(clock), .in1(R8375));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8541 (.out1(R8542), .clock(clock), .in1(R8541));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8702 (.out1(R8703), .clock(clock), .in1(R8702));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8910 (.out1(R8911), .clock(clock), .in1(R8910));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9063 (.out1(R9064), .clock(clock), .in1(R9063));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9211 (.out1(R9212), .clock(clock), .in1(R9211));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9406 (.out1(R9407), .clock(clock), .in1(R9406));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9546 (.out1(R9547), .clock(clock), .in1(R9546));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9681 (.out1(R9682), .clock(clock), .in1(R9681));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9863 (.out1(R9864), .clock(clock), .in1(R9863));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9990 (.out1(R9991), .clock(clock), .in1(R9990));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10112 (.out1(R10113), .clock(clock), .in1(R10112));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10281 (.out1(R10282), .clock(clock), .in1(R10281));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10394 (.out1(R10395), .clock(clock), .in1(R10394));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10502 (.out1(R10503), .clock(clock), .in1(R10502));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10643 (.out1(R10644), .clock(clock), .in1(_1013));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10644 (.out1(R10645), .clock(clock), .in1(_993));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10645 (.out1(R10646), .clock(clock), .in1(_982));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10646 (.out1(R10647), .clock(clock), .in1(_975));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10647 (.out1(R10648), .clock(clock), .in1(_976));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10648 (.out1(R10649), .clock(clock), .in1(_1044));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10649 (.out1(R10650), .clock(clock), .in1(_1024));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10650 (.out1(R10651), .clock(clock), .in1(_1015));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10651 (.out1(R10652), .clock(clock), .in1(_1004));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10652 (.out1(R10653), .clock(clock), .in1(_995));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10653 (.out1(R10654), .clock(clock), .in1(_984));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1059 (.out1(_1025), .in1(R10650), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1050 (.out1(_1016), .in1(R10644), .in2(R10651));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1019 (.out1(_985), .in1(R10646), .in2(R10654));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1079 (.out1(_1045), .in1(R10649), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1060 (.out1(_1026), .in1(_1016), .in2(_1025));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1039 (.out1(_1005), .in1(R10652), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1030 (.out1(_996), .in1(R10645), .in2(R10653));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1020 (.out1(_986), .in1(_985), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1011 (.out1(_977), .in1(R10648), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1040 (.out1(_1006), .in1(_996), .in2(_1005));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1080 (.out1(_1046), .in1(_1045), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1061 (.out1(_1027), .in1(_1026), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1021 (.out1(_987), .in1(_986), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1012 (.out1(_978), .in1(R10647), .in2(_977));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1081 (.out1(_1047), .in1(_1027), .in2(_1046));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1041 (.out1(_1007), .in1(_1006), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1022 (.out1(_988), .in1(_978), .in2(_987));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3829 (.out1(R3830), .clock(clock), .in1(R3829));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4085 (.out1(R4086), .clock(clock), .in1(R4085));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4340 (.out1(R4341), .clock(clock), .in1(R4340));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4585 (.out1(R4586), .clock(clock), .in1(R4585));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4825 (.out1(R4826), .clock(clock), .in1(R4825));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5112 (.out1(R5113), .clock(clock), .in1(R5112));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5344 (.out1(R5345), .clock(clock), .in1(R5344));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5571 (.out1(R5572), .clock(clock), .in1(R5571));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5845 (.out1(R5846), .clock(clock), .in1(R5845));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6063 (.out1(R6064), .clock(clock), .in1(R6063));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6276 (.out1(R6277), .clock(clock), .in1(R6276));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6537 (.out1(R6538), .clock(clock), .in1(R6537));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6742 (.out1(R6743), .clock(clock), .in1(R6742));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6942 (.out1(R6943), .clock(clock), .in1(R6942));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7189 (.out1(R7190), .clock(clock), .in1(R7189));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7381 (.out1(R7382), .clock(clock), .in1(R7381));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7568 (.out1(R7569), .clock(clock), .in1(R7568));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7802 (.out1(R7803), .clock(clock), .in1(R7802));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7981 (.out1(R7982), .clock(clock), .in1(R7981));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8155 (.out1(R8156), .clock(clock), .in1(R8155));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8376 (.out1(R8377), .clock(clock), .in1(R8376));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8542 (.out1(R8543), .clock(clock), .in1(R8542));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8703 (.out1(R8704), .clock(clock), .in1(R8703));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8911 (.out1(R8912), .clock(clock), .in1(R8911));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9064 (.out1(R9065), .clock(clock), .in1(R9064));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9212 (.out1(R9213), .clock(clock), .in1(R9212));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9407 (.out1(R9408), .clock(clock), .in1(R9407));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9547 (.out1(R9548), .clock(clock), .in1(R9547));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9682 (.out1(R9683), .clock(clock), .in1(R9682));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9864 (.out1(R9865), .clock(clock), .in1(R9864));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9991 (.out1(R9992), .clock(clock), .in1(R9991));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10113 (.out1(R10114), .clock(clock), .in1(R10113));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10282 (.out1(R10283), .clock(clock), .in1(R10282));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10395 (.out1(R10396), .clock(clock), .in1(R10395));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10503 (.out1(R10504), .clock(clock), .in1(R10503));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10654 (.out1(R10655), .clock(clock), .in1(_1047));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10655 (.out1(R10656), .clock(clock), .in1(_1007));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10656 (.out1(R10657), .clock(clock), .in1(_988));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1002 (.out1(_968), .in1(R10283));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1042 (.out1(_1008), .in1(R10656), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1023 (.out1(_989), .in1(R10657), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op1082 (.out1(_1048), .in1(R10655), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1043 (.out1(_1009), .in1(_989), .in2(_1008));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1003 (.out1(_969), .in1(_968), .in2(2 'd 2));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1083 (.out1(_1049), .in1(_1009), .in2(_1048));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op1084 (.out1(_1050), .in1(_1049), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3830 (.out1(R3831), .clock(clock), .in1(R3830));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4086 (.out1(R4087), .clock(clock), .in1(R4086));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4341 (.out1(R4342), .clock(clock), .in1(R4341));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4586 (.out1(R4587), .clock(clock), .in1(R4586));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4826 (.out1(R4827), .clock(clock), .in1(R4826));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5113 (.out1(R5114), .clock(clock), .in1(R5113));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5345 (.out1(R5346), .clock(clock), .in1(R5345));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5572 (.out1(R5573), .clock(clock), .in1(R5572));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5846 (.out1(R5847), .clock(clock), .in1(R5846));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6064 (.out1(R6065), .clock(clock), .in1(R6064));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6277 (.out1(R6278), .clock(clock), .in1(R6277));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6538 (.out1(R6539), .clock(clock), .in1(R6538));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6743 (.out1(R6744), .clock(clock), .in1(R6743));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6943 (.out1(R6944), .clock(clock), .in1(R6943));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7190 (.out1(R7191), .clock(clock), .in1(R7190));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7382 (.out1(R7383), .clock(clock), .in1(R7382));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7569 (.out1(R7570), .clock(clock), .in1(R7569));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7803 (.out1(R7804), .clock(clock), .in1(R7803));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7982 (.out1(R7983), .clock(clock), .in1(R7982));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8156 (.out1(R8157), .clock(clock), .in1(R8156));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8377 (.out1(R8378), .clock(clock), .in1(R8377));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8543 (.out1(R8544), .clock(clock), .in1(R8543));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8704 (.out1(R8705), .clock(clock), .in1(R8704));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8912 (.out1(R8913), .clock(clock), .in1(R8912));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9065 (.out1(R9066), .clock(clock), .in1(R9065));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9213 (.out1(R9214), .clock(clock), .in1(R9213));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9408 (.out1(R9409), .clock(clock), .in1(R9408));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9548 (.out1(R9549), .clock(clock), .in1(R9548));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9683 (.out1(R9684), .clock(clock), .in1(R9683));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9865 (.out1(R9866), .clock(clock), .in1(R9865));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9992 (.out1(R9993), .clock(clock), .in1(R9992));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10114 (.out1(R10115), .clock(clock), .in1(R10114));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10283 (.out1(R10284), .clock(clock), .in1(R10283));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10396 (.out1(R10397), .clock(clock), .in1(R10396));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10504 (.out1(R10505), .clock(clock), .in1(R10504));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10657 (.out1(R10658), .clock(clock), .in1(_969));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10658 (.out1(R10659), .clock(clock), .in1(_1050));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op1085 (.out1(_1051), .in1(R10659), .in2(57 'd 72340172838076673));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1004 (.out1(_970), .in1(base0_76_3625_D), .in2(R10658));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3831 (.out1(R3832), .clock(clock), .in1(R3831));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4087 (.out1(R4088), .clock(clock), .in1(R4087));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4342 (.out1(R4343), .clock(clock), .in1(R4342));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4587 (.out1(R4588), .clock(clock), .in1(R4587));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4827 (.out1(R4828), .clock(clock), .in1(R4827));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5114 (.out1(R5115), .clock(clock), .in1(R5114));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5346 (.out1(R5347), .clock(clock), .in1(R5346));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5573 (.out1(R5574), .clock(clock), .in1(R5573));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5847 (.out1(R5848), .clock(clock), .in1(R5847));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6065 (.out1(R6066), .clock(clock), .in1(R6065));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6278 (.out1(R6279), .clock(clock), .in1(R6278));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6539 (.out1(R6540), .clock(clock), .in1(R6539));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6744 (.out1(R6745), .clock(clock), .in1(R6744));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6944 (.out1(R6945), .clock(clock), .in1(R6944));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7191 (.out1(R7192), .clock(clock), .in1(R7191));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7383 (.out1(R7384), .clock(clock), .in1(R7383));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7570 (.out1(R7571), .clock(clock), .in1(R7570));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7804 (.out1(R7805), .clock(clock), .in1(R7804));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7983 (.out1(R7984), .clock(clock), .in1(R7983));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8157 (.out1(R8158), .clock(clock), .in1(R8157));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8378 (.out1(R8379), .clock(clock), .in1(R8378));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8544 (.out1(R8545), .clock(clock), .in1(R8544));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8705 (.out1(R8706), .clock(clock), .in1(R8705));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8913 (.out1(R8914), .clock(clock), .in1(R8913));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9066 (.out1(R9067), .clock(clock), .in1(R9066));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9214 (.out1(R9215), .clock(clock), .in1(R9214));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9409 (.out1(R9410), .clock(clock), .in1(R9409));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9549 (.out1(R9550), .clock(clock), .in1(R9549));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9684 (.out1(R9685), .clock(clock), .in1(R9684));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9866 (.out1(R9867), .clock(clock), .in1(R9866));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9993 (.out1(R9994), .clock(clock), .in1(R9993));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10115 (.out1(R10116), .clock(clock), .in1(R10115));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10284 (.out1(R10285), .clock(clock), .in1(R10284));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10397 (.out1(R10398), .clock(clock), .in1(R10397));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10505 (.out1(R10506), .clock(clock), .in1(R10505));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10659 (.out1(R10660), .clock(clock), .in1(_1051));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10660 (.out1(R10661), .clock(clock), .in1(_970));
  SRAM op1005 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_971),.ADR(R10661));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op1086 (.out1(_1052), .in1(R10660), .in2(6 'd 56));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3832 (.out1(R3833), .clock(clock), .in1(R3832));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4088 (.out1(R4089), .clock(clock), .in1(R4088));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4343 (.out1(R4344), .clock(clock), .in1(R4343));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4588 (.out1(R4589), .clock(clock), .in1(R4588));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4828 (.out1(R4829), .clock(clock), .in1(R4828));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5115 (.out1(R5116), .clock(clock), .in1(R5115));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5347 (.out1(R5348), .clock(clock), .in1(R5347));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5574 (.out1(R5575), .clock(clock), .in1(R5574));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5848 (.out1(R5849), .clock(clock), .in1(R5848));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6066 (.out1(R6067), .clock(clock), .in1(R6066));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6279 (.out1(R6280), .clock(clock), .in1(R6279));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6540 (.out1(R6541), .clock(clock), .in1(R6540));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6745 (.out1(R6746), .clock(clock), .in1(R6745));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6945 (.out1(R6946), .clock(clock), .in1(R6945));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7192 (.out1(R7193), .clock(clock), .in1(R7192));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7384 (.out1(R7385), .clock(clock), .in1(R7384));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7571 (.out1(R7572), .clock(clock), .in1(R7571));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7805 (.out1(R7806), .clock(clock), .in1(R7805));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7984 (.out1(R7985), .clock(clock), .in1(R7984));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8158 (.out1(R8159), .clock(clock), .in1(R8158));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8379 (.out1(R8380), .clock(clock), .in1(R8379));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8545 (.out1(R8546), .clock(clock), .in1(R8545));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8706 (.out1(R8707), .clock(clock), .in1(R8706));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8914 (.out1(R8915), .clock(clock), .in1(R8914));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9067 (.out1(R9068), .clock(clock), .in1(R9067));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9215 (.out1(R9216), .clock(clock), .in1(R9215));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9410 (.out1(R9411), .clock(clock), .in1(R9410));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9550 (.out1(R9551), .clock(clock), .in1(R9550));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9685 (.out1(R9686), .clock(clock), .in1(R9685));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9867 (.out1(R9868), .clock(clock), .in1(R9867));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9994 (.out1(R9995), .clock(clock), .in1(R9994));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10116 (.out1(R10117), .clock(clock), .in1(R10116));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10285 (.out1(R10286), .clock(clock), .in1(R10285));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10398 (.out1(R10399), .clock(clock), .in1(R10398));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10506 (.out1(R10507), .clock(clock), .in1(R10506));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10661 (.out1(R10662), .clock(clock), .in1(_971));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10662 (.out1(R10663), .clock(clock), .in1(_1052));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1087 (.out1(_1053), .in1(R10663));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1088 (.out1(_1054), .in1(R10662), .in2(_1053));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1089 (.out1(idx_3626), .in1(_1054), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3833 (.out1(R3834), .clock(clock), .in1(R3833));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4089 (.out1(R4090), .clock(clock), .in1(R4089));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4344 (.out1(R4345), .clock(clock), .in1(R4344));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4589 (.out1(R4590), .clock(clock), .in1(R4589));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4829 (.out1(R4830), .clock(clock), .in1(R4829));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5116 (.out1(R5117), .clock(clock), .in1(R5116));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5348 (.out1(R5349), .clock(clock), .in1(R5348));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5575 (.out1(R5576), .clock(clock), .in1(R5575));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5849 (.out1(R5850), .clock(clock), .in1(R5849));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6067 (.out1(R6068), .clock(clock), .in1(R6067));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6280 (.out1(R6281), .clock(clock), .in1(R6280));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6541 (.out1(R6542), .clock(clock), .in1(R6541));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6746 (.out1(R6747), .clock(clock), .in1(R6746));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6946 (.out1(R6947), .clock(clock), .in1(R6946));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7193 (.out1(R7194), .clock(clock), .in1(R7193));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7385 (.out1(R7386), .clock(clock), .in1(R7385));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7572 (.out1(R7573), .clock(clock), .in1(R7572));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7806 (.out1(R7807), .clock(clock), .in1(R7806));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7985 (.out1(R7986), .clock(clock), .in1(R7985));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8159 (.out1(R8160), .clock(clock), .in1(R8159));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8380 (.out1(R8381), .clock(clock), .in1(R8380));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8546 (.out1(R8547), .clock(clock), .in1(R8546));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8707 (.out1(R8708), .clock(clock), .in1(R8707));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8915 (.out1(R8916), .clock(clock), .in1(R8915));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9068 (.out1(R9069), .clock(clock), .in1(R9068));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9216 (.out1(R9217), .clock(clock), .in1(R9216));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9411 (.out1(R9412), .clock(clock), .in1(R9411));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9551 (.out1(R9552), .clock(clock), .in1(R9551));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9686 (.out1(R9687), .clock(clock), .in1(R9686));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9868 (.out1(R9869), .clock(clock), .in1(R9868));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9995 (.out1(R9996), .clock(clock), .in1(R9995));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10117 (.out1(R10118), .clock(clock), .in1(R10117));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10286 (.out1(R10287), .clock(clock), .in1(R10286));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10399 (.out1(R10400), .clock(clock), .in1(R10399));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10507 (.out1(R10508), .clock(clock), .in1(R10507));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10663 (.out1(R10664), .clock(clock), .in1(idx_3626));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1093 (.out1(_1057), .in1(R10664));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1094 (.out1(_1058), .in1(_1057), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3834 (.out1(R3835), .clock(clock), .in1(R3834));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4090 (.out1(R4091), .clock(clock), .in1(R4090));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4345 (.out1(R4346), .clock(clock), .in1(R4345));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4590 (.out1(R4591), .clock(clock), .in1(R4590));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4830 (.out1(R4831), .clock(clock), .in1(R4830));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5117 (.out1(R5118), .clock(clock), .in1(R5117));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5349 (.out1(R5350), .clock(clock), .in1(R5349));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5576 (.out1(R5577), .clock(clock), .in1(R5576));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5850 (.out1(R5851), .clock(clock), .in1(R5850));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6068 (.out1(R6069), .clock(clock), .in1(R6068));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6281 (.out1(R6282), .clock(clock), .in1(R6281));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6542 (.out1(R6543), .clock(clock), .in1(R6542));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6747 (.out1(R6748), .clock(clock), .in1(R6747));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6947 (.out1(R6948), .clock(clock), .in1(R6947));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7194 (.out1(R7195), .clock(clock), .in1(R7194));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7386 (.out1(R7387), .clock(clock), .in1(R7386));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7573 (.out1(R7574), .clock(clock), .in1(R7573));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7807 (.out1(R7808), .clock(clock), .in1(R7807));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7986 (.out1(R7987), .clock(clock), .in1(R7986));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8160 (.out1(R8161), .clock(clock), .in1(R8160));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8381 (.out1(R8382), .clock(clock), .in1(R8381));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8547 (.out1(R8548), .clock(clock), .in1(R8547));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8708 (.out1(R8709), .clock(clock), .in1(R8708));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8916 (.out1(R8917), .clock(clock), .in1(R8916));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9069 (.out1(R9070), .clock(clock), .in1(R9069));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9217 (.out1(R9218), .clock(clock), .in1(R9217));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9412 (.out1(R9413), .clock(clock), .in1(R9412));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9552 (.out1(R9553), .clock(clock), .in1(R9552));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9687 (.out1(R9688), .clock(clock), .in1(R9687));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9869 (.out1(R9870), .clock(clock), .in1(R9869));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9996 (.out1(R9997), .clock(clock), .in1(R9996));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10118 (.out1(R10119), .clock(clock), .in1(R10118));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10287 (.out1(R10288), .clock(clock), .in1(R10287));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10400 (.out1(R10401), .clock(clock), .in1(R10400));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10508 (.out1(R10509), .clock(clock), .in1(R10508));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10664 (.out1(R10665), .clock(clock), .in1(R10664));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10764 (.out1(R10765), .clock(clock), .in1(_1058));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1095 (.out1(_1059), .in1(vec82_3628_D), .in2(R10765));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3835 (.out1(R3836), .clock(clock), .in1(R3835));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4091 (.out1(R4092), .clock(clock), .in1(R4091));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4346 (.out1(R4347), .clock(clock), .in1(R4346));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4591 (.out1(R4592), .clock(clock), .in1(R4591));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4831 (.out1(R4832), .clock(clock), .in1(R4831));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5118 (.out1(R5119), .clock(clock), .in1(R5118));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5350 (.out1(R5351), .clock(clock), .in1(R5350));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5577 (.out1(R5578), .clock(clock), .in1(R5577));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5851 (.out1(R5852), .clock(clock), .in1(R5851));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6069 (.out1(R6070), .clock(clock), .in1(R6069));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6282 (.out1(R6283), .clock(clock), .in1(R6282));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6543 (.out1(R6544), .clock(clock), .in1(R6543));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6748 (.out1(R6749), .clock(clock), .in1(R6748));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6948 (.out1(R6949), .clock(clock), .in1(R6948));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7195 (.out1(R7196), .clock(clock), .in1(R7195));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7387 (.out1(R7388), .clock(clock), .in1(R7387));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7574 (.out1(R7575), .clock(clock), .in1(R7574));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7808 (.out1(R7809), .clock(clock), .in1(R7808));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7987 (.out1(R7988), .clock(clock), .in1(R7987));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8161 (.out1(R8162), .clock(clock), .in1(R8161));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8382 (.out1(R8383), .clock(clock), .in1(R8382));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8548 (.out1(R8549), .clock(clock), .in1(R8548));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8709 (.out1(R8710), .clock(clock), .in1(R8709));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8917 (.out1(R8918), .clock(clock), .in1(R8917));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9070 (.out1(R9071), .clock(clock), .in1(R9070));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9218 (.out1(R9219), .clock(clock), .in1(R9218));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9413 (.out1(R9414), .clock(clock), .in1(R9413));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9553 (.out1(R9554), .clock(clock), .in1(R9553));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9688 (.out1(R9689), .clock(clock), .in1(R9688));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9870 (.out1(R9871), .clock(clock), .in1(R9870));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9997 (.out1(R9998), .clock(clock), .in1(R9997));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10119 (.out1(R10120), .clock(clock), .in1(R10119));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10288 (.out1(R10289), .clock(clock), .in1(R10288));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10401 (.out1(R10402), .clock(clock), .in1(R10401));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10509 (.out1(R10510), .clock(clock), .in1(R10509));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10665 (.out1(R10666), .clock(clock), .in1(R10665));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10765 (.out1(R10766), .clock(clock), .in1(_1059));
  SRAM op1096 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1060),.ADR(R10766));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3836 (.out1(R3837), .clock(clock), .in1(R3836));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4092 (.out1(R4093), .clock(clock), .in1(R4092));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4347 (.out1(R4348), .clock(clock), .in1(R4347));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4592 (.out1(R4593), .clock(clock), .in1(R4592));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4832 (.out1(R4833), .clock(clock), .in1(R4832));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5119 (.out1(R5120), .clock(clock), .in1(R5119));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5351 (.out1(R5352), .clock(clock), .in1(R5351));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5578 (.out1(R5579), .clock(clock), .in1(R5578));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5852 (.out1(R5853), .clock(clock), .in1(R5852));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6070 (.out1(R6071), .clock(clock), .in1(R6070));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6283 (.out1(R6284), .clock(clock), .in1(R6283));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6544 (.out1(R6545), .clock(clock), .in1(R6544));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6749 (.out1(R6750), .clock(clock), .in1(R6749));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6949 (.out1(R6950), .clock(clock), .in1(R6949));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7196 (.out1(R7197), .clock(clock), .in1(R7196));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7388 (.out1(R7389), .clock(clock), .in1(R7388));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7575 (.out1(R7576), .clock(clock), .in1(R7575));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7809 (.out1(R7810), .clock(clock), .in1(R7809));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7988 (.out1(R7989), .clock(clock), .in1(R7988));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8162 (.out1(R8163), .clock(clock), .in1(R8162));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8383 (.out1(R8384), .clock(clock), .in1(R8383));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8549 (.out1(R8550), .clock(clock), .in1(R8549));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8710 (.out1(R8711), .clock(clock), .in1(R8710));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8918 (.out1(R8919), .clock(clock), .in1(R8918));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9071 (.out1(R9072), .clock(clock), .in1(R9071));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9219 (.out1(R9220), .clock(clock), .in1(R9219));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9414 (.out1(R9415), .clock(clock), .in1(R9414));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9554 (.out1(R9555), .clock(clock), .in1(R9554));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9689 (.out1(R9690), .clock(clock), .in1(R9689));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9871 (.out1(R9872), .clock(clock), .in1(R9871));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9998 (.out1(R9999), .clock(clock), .in1(R9998));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10120 (.out1(R10121), .clock(clock), .in1(R10120));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10289 (.out1(R10290), .clock(clock), .in1(R10289));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10402 (.out1(R10403), .clock(clock), .in1(R10402));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10510 (.out1(R10511), .clock(clock), .in1(R10510));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10666 (.out1(R10667), .clock(clock), .in1(R10666));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10766 (.out1(R10767), .clock(clock), .in1(_1060));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op1090 (.out1(_1055), .in1(ip2_3602_D), .in2(6 'd 40));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1091 (.out1(_1056), .in1(_1055));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op1092 (.out1(off_3627), .in1(_1056), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1097 (.out1(_1061), .in1(R10767), .in2(off_3627));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3837 (.out1(R3838), .clock(clock), .in1(R3837));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4093 (.out1(R4094), .clock(clock), .in1(R4093));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4348 (.out1(R4349), .clock(clock), .in1(R4348));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4593 (.out1(R4594), .clock(clock), .in1(R4593));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4833 (.out1(R4834), .clock(clock), .in1(R4833));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5120 (.out1(R5121), .clock(clock), .in1(R5120));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5352 (.out1(R5353), .clock(clock), .in1(R5352));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5579 (.out1(R5580), .clock(clock), .in1(R5579));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5853 (.out1(R5854), .clock(clock), .in1(R5853));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6071 (.out1(R6072), .clock(clock), .in1(R6071));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6284 (.out1(R6285), .clock(clock), .in1(R6284));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6545 (.out1(R6546), .clock(clock), .in1(R6545));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6750 (.out1(R6751), .clock(clock), .in1(R6750));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6950 (.out1(R6951), .clock(clock), .in1(R6950));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7197 (.out1(R7198), .clock(clock), .in1(R7197));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7389 (.out1(R7390), .clock(clock), .in1(R7389));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7576 (.out1(R7577), .clock(clock), .in1(R7576));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7810 (.out1(R7811), .clock(clock), .in1(R7810));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7989 (.out1(R7990), .clock(clock), .in1(R7989));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8163 (.out1(R8164), .clock(clock), .in1(R8163));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8384 (.out1(R8385), .clock(clock), .in1(R8384));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8550 (.out1(R8551), .clock(clock), .in1(R8550));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8711 (.out1(R8712), .clock(clock), .in1(R8711));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8919 (.out1(R8920), .clock(clock), .in1(R8919));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9072 (.out1(R9073), .clock(clock), .in1(R9072));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9220 (.out1(R9221), .clock(clock), .in1(R9220));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9415 (.out1(R9416), .clock(clock), .in1(R9415));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9555 (.out1(R9556), .clock(clock), .in1(R9555));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9690 (.out1(R9691), .clock(clock), .in1(R9690));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9872 (.out1(R9873), .clock(clock), .in1(R9872));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9999 (.out1(R10000), .clock(clock), .in1(R9999));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10121 (.out1(R10122), .clock(clock), .in1(R10121));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10290 (.out1(R10291), .clock(clock), .in1(R10290));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10403 (.out1(R10404), .clock(clock), .in1(R10403));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10511 (.out1(R10512), .clock(clock), .in1(R10511));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10667 (.out1(R10668), .clock(clock), .in1(R10667));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10767 (.out1(R10768), .clock(clock), .in1(off_3627));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10862 (.out1(R10863), .clock(clock), .in1(_1061));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op1098 (.out1(_1062), .in1(R10863), .in2(1 'd 1));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op1099 (.out1(ifout1099), .in1(_1062), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1167 (.out1(_1130), .in1(R10668));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1160 (.out1(_1123), .in1(R10668));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1149 (.out1(_1112), .in1(R10668));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1129 (.out1(_1092), .in1(R10668));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1168 (.out1(_1131), .in1(_1130), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1161 (.out1(_1124), .in1(_1123), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1150 (.out1(_1113), .in1(_1112), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1130 (.out1(_1093), .in1(_1092), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3838 (.out1(R3839), .clock(clock), .in1(R3838));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4094 (.out1(R4095), .clock(clock), .in1(R4094));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4349 (.out1(R4350), .clock(clock), .in1(R4349));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4594 (.out1(R4595), .clock(clock), .in1(R4594));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4834 (.out1(R4835), .clock(clock), .in1(R4834));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5121 (.out1(R5122), .clock(clock), .in1(R5121));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5353 (.out1(R5354), .clock(clock), .in1(R5353));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5580 (.out1(R5581), .clock(clock), .in1(R5580));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5854 (.out1(R5855), .clock(clock), .in1(R5854));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6072 (.out1(R6073), .clock(clock), .in1(R6072));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6285 (.out1(R6286), .clock(clock), .in1(R6285));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6546 (.out1(R6547), .clock(clock), .in1(R6546));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6751 (.out1(R6752), .clock(clock), .in1(R6751));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6951 (.out1(R6952), .clock(clock), .in1(R6951));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7198 (.out1(R7199), .clock(clock), .in1(R7198));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7390 (.out1(R7391), .clock(clock), .in1(R7390));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7577 (.out1(R7578), .clock(clock), .in1(R7577));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7811 (.out1(R7812), .clock(clock), .in1(R7811));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7990 (.out1(R7991), .clock(clock), .in1(R7990));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8164 (.out1(R8165), .clock(clock), .in1(R8164));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8385 (.out1(R8386), .clock(clock), .in1(R8385));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8551 (.out1(R8552), .clock(clock), .in1(R8551));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8712 (.out1(R8713), .clock(clock), .in1(R8712));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8920 (.out1(R8921), .clock(clock), .in1(R8920));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9073 (.out1(R9074), .clock(clock), .in1(R9073));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9221 (.out1(R9222), .clock(clock), .in1(R9221));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9416 (.out1(R9417), .clock(clock), .in1(R9416));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9556 (.out1(R9557), .clock(clock), .in1(R9556));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9691 (.out1(R9692), .clock(clock), .in1(R9691));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9873 (.out1(R9874), .clock(clock), .in1(R9873));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10000 (.out1(R10001), .clock(clock), .in1(R10000));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10122 (.out1(R10123), .clock(clock), .in1(R10122));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10291 (.out1(R10292), .clock(clock), .in1(R10291));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10404 (.out1(R10405), .clock(clock), .in1(R10404));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10512 (.out1(R10513), .clock(clock), .in1(R10512));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10668 (.out1(R10669), .clock(clock), .in1(R10668));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10768 (.out1(R10769), .clock(clock), .in1(R10768));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10863 (.out1(R10864), .clock(clock), .in1(ifout1099));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10965 (.out1(R10966), .clock(clock), .in1(_1131));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10966 (.out1(R10967), .clock(clock), .in1(_1124));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10967 (.out1(R10968), .clock(clock), .in1(_1113));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10968 (.out1(R10969), .clock(clock), .in1(_1093));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1142 (.out1(_1105), .in1(R10669));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1122 (.out1(_1085), .in1(R10669));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1111 (.out1(_1074), .in1(R10669));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1104 (.out1(_1067), .in1(R10669));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1171 (.out1(_1134), .in1(2 'd 2), .in2(R10769));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1143 (.out1(_1106), .in1(_1105), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1123 (.out1(_1086), .in1(_1085), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1112 (.out1(_1075), .in1(_1074), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1105 (.out1(_1068), .in1(_1067), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1169 (.out1(_1132), .in1(vec82_3628_D), .in2(R10966));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1162 (.out1(_1125), .in1(vec82_3628_D), .in2(R10967));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1151 (.out1(_1114), .in1(vec82_3628_D), .in2(R10968));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1131 (.out1(_1094), .in1(vec82_3628_D), .in2(R10969));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3839 (.out1(R3840), .clock(clock), .in1(R3839));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4095 (.out1(R4096), .clock(clock), .in1(R4095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4350 (.out1(R4351), .clock(clock), .in1(R4350));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4595 (.out1(R4596), .clock(clock), .in1(R4595));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4835 (.out1(R4836), .clock(clock), .in1(R4835));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5122 (.out1(R5123), .clock(clock), .in1(R5122));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5354 (.out1(R5355), .clock(clock), .in1(R5354));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5581 (.out1(R5582), .clock(clock), .in1(R5581));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5855 (.out1(R5856), .clock(clock), .in1(R5855));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6073 (.out1(R6074), .clock(clock), .in1(R6073));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6286 (.out1(R6287), .clock(clock), .in1(R6286));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6547 (.out1(R6548), .clock(clock), .in1(R6547));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6752 (.out1(R6753), .clock(clock), .in1(R6752));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6952 (.out1(R6953), .clock(clock), .in1(R6952));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7199 (.out1(R7200), .clock(clock), .in1(R7199));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7391 (.out1(R7392), .clock(clock), .in1(R7391));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7578 (.out1(R7579), .clock(clock), .in1(R7578));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7812 (.out1(R7813), .clock(clock), .in1(R7812));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7991 (.out1(R7992), .clock(clock), .in1(R7991));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8165 (.out1(R8166), .clock(clock), .in1(R8165));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8386 (.out1(R8387), .clock(clock), .in1(R8386));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8552 (.out1(R8553), .clock(clock), .in1(R8552));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8713 (.out1(R8714), .clock(clock), .in1(R8713));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8921 (.out1(R8922), .clock(clock), .in1(R8921));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9074 (.out1(R9075), .clock(clock), .in1(R9074));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9222 (.out1(R9223), .clock(clock), .in1(R9222));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9417 (.out1(R9418), .clock(clock), .in1(R9417));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9557 (.out1(R9558), .clock(clock), .in1(R9557));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9692 (.out1(R9693), .clock(clock), .in1(R9692));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9874 (.out1(R9875), .clock(clock), .in1(R9874));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10001 (.out1(R10002), .clock(clock), .in1(R10001));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10123 (.out1(R10124), .clock(clock), .in1(R10123));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10292 (.out1(R10293), .clock(clock), .in1(R10292));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10405 (.out1(R10406), .clock(clock), .in1(R10405));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10513 (.out1(R10514), .clock(clock), .in1(R10513));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10669 (.out1(R10670), .clock(clock), .in1(R10669));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10769 (.out1(R10770), .clock(clock), .in1(R10769));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10864 (.out1(R10865), .clock(clock), .in1(R10864));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10969 (.out1(R10970), .clock(clock), .in1(_1134));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10970 (.out1(R10971), .clock(clock), .in1(_1106));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10971 (.out1(R10972), .clock(clock), .in1(_1086));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10972 (.out1(R10973), .clock(clock), .in1(_1075));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10973 (.out1(R10974), .clock(clock), .in1(_1068));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10974 (.out1(R10975), .clock(clock), .in1(_1132));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10975 (.out1(R10976), .clock(clock), .in1(_1125));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10976 (.out1(R10977), .clock(clock), .in1(_1114));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10977 (.out1(R10978), .clock(clock), .in1(_1094));
  SRAM op1170 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1133),.ADR(R10975));
  SRAM op1163 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1126),.ADR(R10976));
  SRAM op1152 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1115),.ADR(R10977));
  SRAM op1132 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1095),.ADR(R10978));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1164 (.out1(_1127), .in1(2 'd 2), .in2(R10770));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1153 (.out1(_1116), .in1(2 'd 2), .in2(R10770));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1146 (.out1(_1109), .in1(2 'd 2), .in2(R10770));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1133 (.out1(_1096), .in1(2 'd 2), .in2(R10770));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1126 (.out1(_1089), .in1(2 'd 2), .in2(R10770));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1115 (.out1(_1078), .in1(2 'd 2), .in2(R10770));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1144 (.out1(_1107), .in1(vec82_3628_D), .in2(R10971));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1124 (.out1(_1087), .in1(vec82_3628_D), .in2(R10972));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1113 (.out1(_1076), .in1(vec82_3628_D), .in2(R10973));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1106 (.out1(_1069), .in1(vec82_3628_D), .in2(R10974));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1172 (.out1(_1135), .in1(R10970), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3840 (.out1(R3841), .clock(clock), .in1(R3840));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4096 (.out1(R4097), .clock(clock), .in1(R4096));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4351 (.out1(R4352), .clock(clock), .in1(R4351));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4596 (.out1(R4597), .clock(clock), .in1(R4596));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4836 (.out1(R4837), .clock(clock), .in1(R4836));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5123 (.out1(R5124), .clock(clock), .in1(R5123));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5355 (.out1(R5356), .clock(clock), .in1(R5355));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5582 (.out1(R5583), .clock(clock), .in1(R5582));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5856 (.out1(R5857), .clock(clock), .in1(R5856));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6074 (.out1(R6075), .clock(clock), .in1(R6074));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6287 (.out1(R6288), .clock(clock), .in1(R6287));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6548 (.out1(R6549), .clock(clock), .in1(R6548));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6753 (.out1(R6754), .clock(clock), .in1(R6753));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6953 (.out1(R6954), .clock(clock), .in1(R6953));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7200 (.out1(R7201), .clock(clock), .in1(R7200));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7392 (.out1(R7393), .clock(clock), .in1(R7392));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7579 (.out1(R7580), .clock(clock), .in1(R7579));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7813 (.out1(R7814), .clock(clock), .in1(R7813));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7992 (.out1(R7993), .clock(clock), .in1(R7992));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8166 (.out1(R8167), .clock(clock), .in1(R8166));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8387 (.out1(R8388), .clock(clock), .in1(R8387));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8553 (.out1(R8554), .clock(clock), .in1(R8553));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8714 (.out1(R8715), .clock(clock), .in1(R8714));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8922 (.out1(R8923), .clock(clock), .in1(R8922));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9075 (.out1(R9076), .clock(clock), .in1(R9075));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9223 (.out1(R9224), .clock(clock), .in1(R9223));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9418 (.out1(R9419), .clock(clock), .in1(R9418));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9558 (.out1(R9559), .clock(clock), .in1(R9558));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9693 (.out1(R9694), .clock(clock), .in1(R9693));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9875 (.out1(R9876), .clock(clock), .in1(R9875));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10002 (.out1(R10003), .clock(clock), .in1(R10002));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10124 (.out1(R10125), .clock(clock), .in1(R10124));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10293 (.out1(R10294), .clock(clock), .in1(R10293));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10406 (.out1(R10407), .clock(clock), .in1(R10406));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10514 (.out1(R10515), .clock(clock), .in1(R10514));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10670 (.out1(R10671), .clock(clock), .in1(R10670));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10770 (.out1(R10771), .clock(clock), .in1(R10770));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10865 (.out1(R10866), .clock(clock), .in1(R10865));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10978 (.out1(R10979), .clock(clock), .in1(_1133));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10979 (.out1(R10980), .clock(clock), .in1(_1126));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10980 (.out1(R10981), .clock(clock), .in1(_1115));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10981 (.out1(R10982), .clock(clock), .in1(_1095));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10982 (.out1(R10983), .clock(clock), .in1(_1127));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10983 (.out1(R10984), .clock(clock), .in1(_1116));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10984 (.out1(R10985), .clock(clock), .in1(_1109));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10985 (.out1(R10986), .clock(clock), .in1(_1096));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10986 (.out1(R10987), .clock(clock), .in1(_1089));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10987 (.out1(R10988), .clock(clock), .in1(_1078));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10988 (.out1(R10989), .clock(clock), .in1(_1107));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10989 (.out1(R10990), .clock(clock), .in1(_1087));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10990 (.out1(R10991), .clock(clock), .in1(_1076));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10991 (.out1(R10992), .clock(clock), .in1(_1069));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10992 (.out1(R10993), .clock(clock), .in1(_1135));
  SRAM op1145 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1108),.ADR(R10989));
  SRAM op1125 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1088),.ADR(R10990));
  SRAM op1114 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1077),.ADR(R10991));
  SRAM op1107 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1070),.ADR(R10992));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1173 (.out1(_1136), .in1(R10979), .in2(R10993));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1174 (.out1(_1137), .in1(_1136), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1165 (.out1(_1128), .in1(R10983), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1154 (.out1(_1117), .in1(R10984), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1134 (.out1(_1097), .in1(R10986), .in2(64 'd 18446744073709551615));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1108 (.out1(_1071), .in1(2 'd 2), .in2(R10771));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1175 (.out1(_1138), .in1(_1137), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1166 (.out1(_1129), .in1(R10980), .in2(_1128));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1155 (.out1(_1118), .in1(R10981), .in2(_1117));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1135 (.out1(_1098), .in1(R10982), .in2(_1097));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1176 (.out1(_1139), .in1(_1129), .in2(_1138));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1156 (.out1(_1119), .in1(_1118), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1147 (.out1(_1110), .in1(R10985), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1136 (.out1(_1099), .in1(_1098), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1127 (.out1(_1090), .in1(R10987), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1116 (.out1(_1079), .in1(R10988), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3841 (.out1(R3842), .clock(clock), .in1(R3841));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4097 (.out1(R4098), .clock(clock), .in1(R4097));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4352 (.out1(R4353), .clock(clock), .in1(R4352));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4597 (.out1(R4598), .clock(clock), .in1(R4597));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4837 (.out1(R4838), .clock(clock), .in1(R4837));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5124 (.out1(R5125), .clock(clock), .in1(R5124));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5356 (.out1(R5357), .clock(clock), .in1(R5356));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5583 (.out1(R5584), .clock(clock), .in1(R5583));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5857 (.out1(R5858), .clock(clock), .in1(R5857));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6075 (.out1(R6076), .clock(clock), .in1(R6075));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6288 (.out1(R6289), .clock(clock), .in1(R6288));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6549 (.out1(R6550), .clock(clock), .in1(R6549));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6754 (.out1(R6755), .clock(clock), .in1(R6754));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6954 (.out1(R6955), .clock(clock), .in1(R6954));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7201 (.out1(R7202), .clock(clock), .in1(R7201));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7393 (.out1(R7394), .clock(clock), .in1(R7393));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7580 (.out1(R7581), .clock(clock), .in1(R7580));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7814 (.out1(R7815), .clock(clock), .in1(R7814));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7993 (.out1(R7994), .clock(clock), .in1(R7993));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8167 (.out1(R8168), .clock(clock), .in1(R8167));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8388 (.out1(R8389), .clock(clock), .in1(R8388));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8554 (.out1(R8555), .clock(clock), .in1(R8554));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8715 (.out1(R8716), .clock(clock), .in1(R8715));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8923 (.out1(R8924), .clock(clock), .in1(R8923));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9076 (.out1(R9077), .clock(clock), .in1(R9076));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9224 (.out1(R9225), .clock(clock), .in1(R9224));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9419 (.out1(R9420), .clock(clock), .in1(R9419));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9559 (.out1(R9560), .clock(clock), .in1(R9559));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9694 (.out1(R9695), .clock(clock), .in1(R9694));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9876 (.out1(R9877), .clock(clock), .in1(R9876));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10003 (.out1(R10004), .clock(clock), .in1(R10003));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10125 (.out1(R10126), .clock(clock), .in1(R10125));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10294 (.out1(R10295), .clock(clock), .in1(R10294));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10407 (.out1(R10408), .clock(clock), .in1(R10407));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10515 (.out1(R10516), .clock(clock), .in1(R10515));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10671 (.out1(R10672), .clock(clock), .in1(R10671));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10771 (.out1(R10772), .clock(clock), .in1(R10771));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10866 (.out1(R10867), .clock(clock), .in1(R10866));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10993 (.out1(R10994), .clock(clock), .in1(_1108));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10994 (.out1(R10995), .clock(clock), .in1(_1088));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10995 (.out1(R10996), .clock(clock), .in1(_1077));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10996 (.out1(R10997), .clock(clock), .in1(_1070));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10997 (.out1(R10998), .clock(clock), .in1(_1071));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10998 (.out1(R10999), .clock(clock), .in1(_1139));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op10999 (.out1(R11000), .clock(clock), .in1(_1119));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11000 (.out1(R11001), .clock(clock), .in1(_1110));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11001 (.out1(R11002), .clock(clock), .in1(_1099));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11002 (.out1(R11003), .clock(clock), .in1(_1090));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11003 (.out1(R11004), .clock(clock), .in1(_1079));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1157 (.out1(_1120), .in1(R11000), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1148 (.out1(_1111), .in1(R10994), .in2(R11001));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1117 (.out1(_1080), .in1(R10996), .in2(R11004));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1177 (.out1(_1140), .in1(R10999), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1158 (.out1(_1121), .in1(_1111), .in2(_1120));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1137 (.out1(_1100), .in1(R11002), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1128 (.out1(_1091), .in1(R10995), .in2(R11003));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1118 (.out1(_1081), .in1(_1080), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1109 (.out1(_1072), .in1(R10998), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1138 (.out1(_1101), .in1(_1091), .in2(_1100));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1178 (.out1(_1141), .in1(_1140), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1159 (.out1(_1122), .in1(_1121), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1119 (.out1(_1082), .in1(_1081), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1110 (.out1(_1073), .in1(R10997), .in2(_1072));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1179 (.out1(_1142), .in1(_1122), .in2(_1141));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1139 (.out1(_1102), .in1(_1101), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1120 (.out1(_1083), .in1(_1073), .in2(_1082));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3842 (.out1(R3843), .clock(clock), .in1(R3842));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4098 (.out1(R4099), .clock(clock), .in1(R4098));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4353 (.out1(R4354), .clock(clock), .in1(R4353));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4598 (.out1(R4599), .clock(clock), .in1(R4598));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4838 (.out1(R4839), .clock(clock), .in1(R4838));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5125 (.out1(R5126), .clock(clock), .in1(R5125));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5357 (.out1(R5358), .clock(clock), .in1(R5357));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5584 (.out1(R5585), .clock(clock), .in1(R5584));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5858 (.out1(R5859), .clock(clock), .in1(R5858));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6076 (.out1(R6077), .clock(clock), .in1(R6076));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6289 (.out1(R6290), .clock(clock), .in1(R6289));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6550 (.out1(R6551), .clock(clock), .in1(R6550));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6755 (.out1(R6756), .clock(clock), .in1(R6755));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6955 (.out1(R6956), .clock(clock), .in1(R6955));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7202 (.out1(R7203), .clock(clock), .in1(R7202));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7394 (.out1(R7395), .clock(clock), .in1(R7394));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7581 (.out1(R7582), .clock(clock), .in1(R7581));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7815 (.out1(R7816), .clock(clock), .in1(R7815));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7994 (.out1(R7995), .clock(clock), .in1(R7994));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8168 (.out1(R8169), .clock(clock), .in1(R8168));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8389 (.out1(R8390), .clock(clock), .in1(R8389));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8555 (.out1(R8556), .clock(clock), .in1(R8555));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8716 (.out1(R8717), .clock(clock), .in1(R8716));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8924 (.out1(R8925), .clock(clock), .in1(R8924));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9077 (.out1(R9078), .clock(clock), .in1(R9077));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9225 (.out1(R9226), .clock(clock), .in1(R9225));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9420 (.out1(R9421), .clock(clock), .in1(R9420));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9560 (.out1(R9561), .clock(clock), .in1(R9560));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9695 (.out1(R9696), .clock(clock), .in1(R9695));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9877 (.out1(R9878), .clock(clock), .in1(R9877));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10004 (.out1(R10005), .clock(clock), .in1(R10004));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10126 (.out1(R10127), .clock(clock), .in1(R10126));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10295 (.out1(R10296), .clock(clock), .in1(R10295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10408 (.out1(R10409), .clock(clock), .in1(R10408));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10516 (.out1(R10517), .clock(clock), .in1(R10516));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10672 (.out1(R10673), .clock(clock), .in1(R10672));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10772 (.out1(R10773), .clock(clock), .in1(R10772));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10867 (.out1(R10868), .clock(clock), .in1(R10867));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11004 (.out1(R11005), .clock(clock), .in1(_1142));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11005 (.out1(R11006), .clock(clock), .in1(_1102));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11006 (.out1(R11007), .clock(clock), .in1(_1083));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1100 (.out1(_1063), .in1(R10673));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1140 (.out1(_1103), .in1(R11006), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1121 (.out1(_1084), .in1(R11007), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op1180 (.out1(_1143), .in1(R11005), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1141 (.out1(_1104), .in1(_1084), .in2(_1103));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1101 (.out1(_1064), .in1(_1063), .in2(2 'd 2));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1181 (.out1(_1144), .in1(_1104), .in2(_1143));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op1182 (.out1(_1145), .in1(_1144), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3843 (.out1(R3844), .clock(clock), .in1(R3843));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4099 (.out1(R4100), .clock(clock), .in1(R4099));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4354 (.out1(R4355), .clock(clock), .in1(R4354));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4599 (.out1(R4600), .clock(clock), .in1(R4599));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4839 (.out1(R4840), .clock(clock), .in1(R4839));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5126 (.out1(R5127), .clock(clock), .in1(R5126));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5358 (.out1(R5359), .clock(clock), .in1(R5358));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5585 (.out1(R5586), .clock(clock), .in1(R5585));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5859 (.out1(R5860), .clock(clock), .in1(R5859));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6077 (.out1(R6078), .clock(clock), .in1(R6077));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6290 (.out1(R6291), .clock(clock), .in1(R6290));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6551 (.out1(R6552), .clock(clock), .in1(R6551));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6756 (.out1(R6757), .clock(clock), .in1(R6756));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6956 (.out1(R6957), .clock(clock), .in1(R6956));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7203 (.out1(R7204), .clock(clock), .in1(R7203));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7395 (.out1(R7396), .clock(clock), .in1(R7395));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7582 (.out1(R7583), .clock(clock), .in1(R7582));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7816 (.out1(R7817), .clock(clock), .in1(R7816));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7995 (.out1(R7996), .clock(clock), .in1(R7995));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8169 (.out1(R8170), .clock(clock), .in1(R8169));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8390 (.out1(R8391), .clock(clock), .in1(R8390));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8556 (.out1(R8557), .clock(clock), .in1(R8556));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8717 (.out1(R8718), .clock(clock), .in1(R8717));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8925 (.out1(R8926), .clock(clock), .in1(R8925));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9078 (.out1(R9079), .clock(clock), .in1(R9078));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9226 (.out1(R9227), .clock(clock), .in1(R9226));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9421 (.out1(R9422), .clock(clock), .in1(R9421));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9561 (.out1(R9562), .clock(clock), .in1(R9561));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9696 (.out1(R9697), .clock(clock), .in1(R9696));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9878 (.out1(R9879), .clock(clock), .in1(R9878));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10005 (.out1(R10006), .clock(clock), .in1(R10005));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10127 (.out1(R10128), .clock(clock), .in1(R10127));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10296 (.out1(R10297), .clock(clock), .in1(R10296));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10409 (.out1(R10410), .clock(clock), .in1(R10409));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10517 (.out1(R10518), .clock(clock), .in1(R10517));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10673 (.out1(R10674), .clock(clock), .in1(R10673));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10773 (.out1(R10774), .clock(clock), .in1(R10773));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10868 (.out1(R10869), .clock(clock), .in1(R10868));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11007 (.out1(R11008), .clock(clock), .in1(_1064));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11008 (.out1(R11009), .clock(clock), .in1(_1145));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op1183 (.out1(_1146), .in1(R11009), .in2(57 'd 72340172838076673));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1102 (.out1(_1065), .in1(base0_82_3633_D), .in2(R11008));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3844 (.out1(R3845), .clock(clock), .in1(R3844));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4100 (.out1(R4101), .clock(clock), .in1(R4100));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4355 (.out1(R4356), .clock(clock), .in1(R4355));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4600 (.out1(R4601), .clock(clock), .in1(R4600));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4840 (.out1(R4841), .clock(clock), .in1(R4840));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5127 (.out1(R5128), .clock(clock), .in1(R5127));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5359 (.out1(R5360), .clock(clock), .in1(R5359));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5586 (.out1(R5587), .clock(clock), .in1(R5586));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5860 (.out1(R5861), .clock(clock), .in1(R5860));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6078 (.out1(R6079), .clock(clock), .in1(R6078));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6291 (.out1(R6292), .clock(clock), .in1(R6291));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6552 (.out1(R6553), .clock(clock), .in1(R6552));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6757 (.out1(R6758), .clock(clock), .in1(R6757));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6957 (.out1(R6958), .clock(clock), .in1(R6957));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7204 (.out1(R7205), .clock(clock), .in1(R7204));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7396 (.out1(R7397), .clock(clock), .in1(R7396));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7583 (.out1(R7584), .clock(clock), .in1(R7583));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7817 (.out1(R7818), .clock(clock), .in1(R7817));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7996 (.out1(R7997), .clock(clock), .in1(R7996));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8170 (.out1(R8171), .clock(clock), .in1(R8170));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8391 (.out1(R8392), .clock(clock), .in1(R8391));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8557 (.out1(R8558), .clock(clock), .in1(R8557));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8718 (.out1(R8719), .clock(clock), .in1(R8718));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8926 (.out1(R8927), .clock(clock), .in1(R8926));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9079 (.out1(R9080), .clock(clock), .in1(R9079));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9227 (.out1(R9228), .clock(clock), .in1(R9227));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9422 (.out1(R9423), .clock(clock), .in1(R9422));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9562 (.out1(R9563), .clock(clock), .in1(R9562));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9697 (.out1(R9698), .clock(clock), .in1(R9697));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9879 (.out1(R9880), .clock(clock), .in1(R9879));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10006 (.out1(R10007), .clock(clock), .in1(R10006));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10128 (.out1(R10129), .clock(clock), .in1(R10128));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10297 (.out1(R10298), .clock(clock), .in1(R10297));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10410 (.out1(R10411), .clock(clock), .in1(R10410));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10518 (.out1(R10519), .clock(clock), .in1(R10518));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10674 (.out1(R10675), .clock(clock), .in1(R10674));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10774 (.out1(R10775), .clock(clock), .in1(R10774));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10869 (.out1(R10870), .clock(clock), .in1(R10869));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11009 (.out1(R11010), .clock(clock), .in1(_1146));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11010 (.out1(R11011), .clock(clock), .in1(_1065));
  SRAM op1103 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1066),.ADR(R11011));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op1184 (.out1(_1147), .in1(R11010), .in2(6 'd 56));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3845 (.out1(R3846), .clock(clock), .in1(R3845));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4101 (.out1(R4102), .clock(clock), .in1(R4101));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4356 (.out1(R4357), .clock(clock), .in1(R4356));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4601 (.out1(R4602), .clock(clock), .in1(R4601));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4841 (.out1(R4842), .clock(clock), .in1(R4841));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5128 (.out1(R5129), .clock(clock), .in1(R5128));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5360 (.out1(R5361), .clock(clock), .in1(R5360));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5587 (.out1(R5588), .clock(clock), .in1(R5587));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5861 (.out1(R5862), .clock(clock), .in1(R5861));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6079 (.out1(R6080), .clock(clock), .in1(R6079));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6292 (.out1(R6293), .clock(clock), .in1(R6292));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6553 (.out1(R6554), .clock(clock), .in1(R6553));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6758 (.out1(R6759), .clock(clock), .in1(R6758));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6958 (.out1(R6959), .clock(clock), .in1(R6958));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7205 (.out1(R7206), .clock(clock), .in1(R7205));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7397 (.out1(R7398), .clock(clock), .in1(R7397));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7584 (.out1(R7585), .clock(clock), .in1(R7584));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7818 (.out1(R7819), .clock(clock), .in1(R7818));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7997 (.out1(R7998), .clock(clock), .in1(R7997));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8171 (.out1(R8172), .clock(clock), .in1(R8171));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8392 (.out1(R8393), .clock(clock), .in1(R8392));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8558 (.out1(R8559), .clock(clock), .in1(R8558));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8719 (.out1(R8720), .clock(clock), .in1(R8719));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8927 (.out1(R8928), .clock(clock), .in1(R8927));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9080 (.out1(R9081), .clock(clock), .in1(R9080));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9228 (.out1(R9229), .clock(clock), .in1(R9228));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9423 (.out1(R9424), .clock(clock), .in1(R9423));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9563 (.out1(R9564), .clock(clock), .in1(R9563));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9698 (.out1(R9699), .clock(clock), .in1(R9698));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9880 (.out1(R9881), .clock(clock), .in1(R9880));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10007 (.out1(R10008), .clock(clock), .in1(R10007));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10129 (.out1(R10130), .clock(clock), .in1(R10129));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10298 (.out1(R10299), .clock(clock), .in1(R10298));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10411 (.out1(R10412), .clock(clock), .in1(R10411));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10519 (.out1(R10520), .clock(clock), .in1(R10519));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10675 (.out1(R10676), .clock(clock), .in1(R10675));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10775 (.out1(R10776), .clock(clock), .in1(R10775));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10870 (.out1(R10871), .clock(clock), .in1(R10870));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11011 (.out1(R11012), .clock(clock), .in1(_1066));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11012 (.out1(R11013), .clock(clock), .in1(_1147));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1185 (.out1(_1148), .in1(R11013));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1186 (.out1(_1149), .in1(R11012), .in2(_1148));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1187 (.out1(idx_3634), .in1(_1149), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3846 (.out1(R3847), .clock(clock), .in1(R3846));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4102 (.out1(R4103), .clock(clock), .in1(R4102));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4357 (.out1(R4358), .clock(clock), .in1(R4357));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4602 (.out1(R4603), .clock(clock), .in1(R4602));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4842 (.out1(R4843), .clock(clock), .in1(R4842));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5129 (.out1(R5130), .clock(clock), .in1(R5129));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5361 (.out1(R5362), .clock(clock), .in1(R5361));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5588 (.out1(R5589), .clock(clock), .in1(R5588));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5862 (.out1(R5863), .clock(clock), .in1(R5862));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6080 (.out1(R6081), .clock(clock), .in1(R6080));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6293 (.out1(R6294), .clock(clock), .in1(R6293));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6554 (.out1(R6555), .clock(clock), .in1(R6554));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6759 (.out1(R6760), .clock(clock), .in1(R6759));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6959 (.out1(R6960), .clock(clock), .in1(R6959));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7206 (.out1(R7207), .clock(clock), .in1(R7206));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7398 (.out1(R7399), .clock(clock), .in1(R7398));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7585 (.out1(R7586), .clock(clock), .in1(R7585));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7819 (.out1(R7820), .clock(clock), .in1(R7819));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7998 (.out1(R7999), .clock(clock), .in1(R7998));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8172 (.out1(R8173), .clock(clock), .in1(R8172));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8393 (.out1(R8394), .clock(clock), .in1(R8393));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8559 (.out1(R8560), .clock(clock), .in1(R8559));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8720 (.out1(R8721), .clock(clock), .in1(R8720));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8928 (.out1(R8929), .clock(clock), .in1(R8928));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9081 (.out1(R9082), .clock(clock), .in1(R9081));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9229 (.out1(R9230), .clock(clock), .in1(R9229));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9424 (.out1(R9425), .clock(clock), .in1(R9424));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9564 (.out1(R9565), .clock(clock), .in1(R9564));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9699 (.out1(R9700), .clock(clock), .in1(R9699));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9881 (.out1(R9882), .clock(clock), .in1(R9881));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10008 (.out1(R10009), .clock(clock), .in1(R10008));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10130 (.out1(R10131), .clock(clock), .in1(R10130));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10299 (.out1(R10300), .clock(clock), .in1(R10299));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10412 (.out1(R10413), .clock(clock), .in1(R10412));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10520 (.out1(R10521), .clock(clock), .in1(R10520));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10676 (.out1(R10677), .clock(clock), .in1(R10676));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10776 (.out1(R10777), .clock(clock), .in1(R10776));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10871 (.out1(R10872), .clock(clock), .in1(R10871));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11013 (.out1(R11014), .clock(clock), .in1(idx_3634));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1191 (.out1(_1152), .in1(R11014));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1192 (.out1(_1153), .in1(_1152), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3847 (.out1(R3848), .clock(clock), .in1(R3847));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4103 (.out1(R4104), .clock(clock), .in1(R4103));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4358 (.out1(R4359), .clock(clock), .in1(R4358));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4603 (.out1(R4604), .clock(clock), .in1(R4603));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4843 (.out1(R4844), .clock(clock), .in1(R4843));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5130 (.out1(R5131), .clock(clock), .in1(R5130));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5362 (.out1(R5363), .clock(clock), .in1(R5362));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5589 (.out1(R5590), .clock(clock), .in1(R5589));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5863 (.out1(R5864), .clock(clock), .in1(R5863));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6081 (.out1(R6082), .clock(clock), .in1(R6081));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6294 (.out1(R6295), .clock(clock), .in1(R6294));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6555 (.out1(R6556), .clock(clock), .in1(R6555));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6760 (.out1(R6761), .clock(clock), .in1(R6760));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6960 (.out1(R6961), .clock(clock), .in1(R6960));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7207 (.out1(R7208), .clock(clock), .in1(R7207));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7399 (.out1(R7400), .clock(clock), .in1(R7399));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7586 (.out1(R7587), .clock(clock), .in1(R7586));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7820 (.out1(R7821), .clock(clock), .in1(R7820));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7999 (.out1(R8000), .clock(clock), .in1(R7999));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8173 (.out1(R8174), .clock(clock), .in1(R8173));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8394 (.out1(R8395), .clock(clock), .in1(R8394));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8560 (.out1(R8561), .clock(clock), .in1(R8560));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8721 (.out1(R8722), .clock(clock), .in1(R8721));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8929 (.out1(R8930), .clock(clock), .in1(R8929));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9082 (.out1(R9083), .clock(clock), .in1(R9082));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9230 (.out1(R9231), .clock(clock), .in1(R9230));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9425 (.out1(R9426), .clock(clock), .in1(R9425));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9565 (.out1(R9566), .clock(clock), .in1(R9565));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9700 (.out1(R9701), .clock(clock), .in1(R9700));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9882 (.out1(R9883), .clock(clock), .in1(R9882));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10009 (.out1(R10010), .clock(clock), .in1(R10009));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10131 (.out1(R10132), .clock(clock), .in1(R10131));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10300 (.out1(R10301), .clock(clock), .in1(R10300));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10413 (.out1(R10414), .clock(clock), .in1(R10413));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10521 (.out1(R10522), .clock(clock), .in1(R10521));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10677 (.out1(R10678), .clock(clock), .in1(R10677));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10777 (.out1(R10778), .clock(clock), .in1(R10777));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10872 (.out1(R10873), .clock(clock), .in1(R10872));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11014 (.out1(R11015), .clock(clock), .in1(R11014));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11101 (.out1(R11102), .clock(clock), .in1(_1153));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1193 (.out1(_1154), .in1(vec88_3636_D), .in2(R11102));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3848 (.out1(R3849), .clock(clock), .in1(R3848));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4104 (.out1(R4105), .clock(clock), .in1(R4104));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4359 (.out1(R4360), .clock(clock), .in1(R4359));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4604 (.out1(R4605), .clock(clock), .in1(R4604));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4844 (.out1(R4845), .clock(clock), .in1(R4844));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5131 (.out1(R5132), .clock(clock), .in1(R5131));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5363 (.out1(R5364), .clock(clock), .in1(R5363));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5590 (.out1(R5591), .clock(clock), .in1(R5590));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5864 (.out1(R5865), .clock(clock), .in1(R5864));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6082 (.out1(R6083), .clock(clock), .in1(R6082));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6295 (.out1(R6296), .clock(clock), .in1(R6295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6556 (.out1(R6557), .clock(clock), .in1(R6556));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6761 (.out1(R6762), .clock(clock), .in1(R6761));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6961 (.out1(R6962), .clock(clock), .in1(R6961));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7208 (.out1(R7209), .clock(clock), .in1(R7208));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7400 (.out1(R7401), .clock(clock), .in1(R7400));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7587 (.out1(R7588), .clock(clock), .in1(R7587));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7821 (.out1(R7822), .clock(clock), .in1(R7821));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8000 (.out1(R8001), .clock(clock), .in1(R8000));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8174 (.out1(R8175), .clock(clock), .in1(R8174));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8395 (.out1(R8396), .clock(clock), .in1(R8395));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8561 (.out1(R8562), .clock(clock), .in1(R8561));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8722 (.out1(R8723), .clock(clock), .in1(R8722));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8930 (.out1(R8931), .clock(clock), .in1(R8930));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9083 (.out1(R9084), .clock(clock), .in1(R9083));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9231 (.out1(R9232), .clock(clock), .in1(R9231));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9426 (.out1(R9427), .clock(clock), .in1(R9426));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9566 (.out1(R9567), .clock(clock), .in1(R9566));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9701 (.out1(R9702), .clock(clock), .in1(R9701));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9883 (.out1(R9884), .clock(clock), .in1(R9883));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10010 (.out1(R10011), .clock(clock), .in1(R10010));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10132 (.out1(R10133), .clock(clock), .in1(R10132));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10301 (.out1(R10302), .clock(clock), .in1(R10301));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10414 (.out1(R10415), .clock(clock), .in1(R10414));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10522 (.out1(R10523), .clock(clock), .in1(R10522));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10678 (.out1(R10679), .clock(clock), .in1(R10678));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10778 (.out1(R10779), .clock(clock), .in1(R10778));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10873 (.out1(R10874), .clock(clock), .in1(R10873));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11015 (.out1(R11016), .clock(clock), .in1(R11015));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11102 (.out1(R11103), .clock(clock), .in1(_1154));
  SRAM op1194 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1155),.ADR(R11103));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3849 (.out1(R3850), .clock(clock), .in1(R3849));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4105 (.out1(R4106), .clock(clock), .in1(R4105));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4360 (.out1(R4361), .clock(clock), .in1(R4360));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4605 (.out1(R4606), .clock(clock), .in1(R4605));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4845 (.out1(R4846), .clock(clock), .in1(R4845));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5132 (.out1(R5133), .clock(clock), .in1(R5132));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5364 (.out1(R5365), .clock(clock), .in1(R5364));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5591 (.out1(R5592), .clock(clock), .in1(R5591));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5865 (.out1(R5866), .clock(clock), .in1(R5865));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6083 (.out1(R6084), .clock(clock), .in1(R6083));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6296 (.out1(R6297), .clock(clock), .in1(R6296));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6557 (.out1(R6558), .clock(clock), .in1(R6557));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6762 (.out1(R6763), .clock(clock), .in1(R6762));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6962 (.out1(R6963), .clock(clock), .in1(R6962));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7209 (.out1(R7210), .clock(clock), .in1(R7209));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7401 (.out1(R7402), .clock(clock), .in1(R7401));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7588 (.out1(R7589), .clock(clock), .in1(R7588));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7822 (.out1(R7823), .clock(clock), .in1(R7822));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8001 (.out1(R8002), .clock(clock), .in1(R8001));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8175 (.out1(R8176), .clock(clock), .in1(R8175));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8396 (.out1(R8397), .clock(clock), .in1(R8396));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8562 (.out1(R8563), .clock(clock), .in1(R8562));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8723 (.out1(R8724), .clock(clock), .in1(R8723));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8931 (.out1(R8932), .clock(clock), .in1(R8931));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9084 (.out1(R9085), .clock(clock), .in1(R9084));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9232 (.out1(R9233), .clock(clock), .in1(R9232));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9427 (.out1(R9428), .clock(clock), .in1(R9427));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9567 (.out1(R9568), .clock(clock), .in1(R9567));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9702 (.out1(R9703), .clock(clock), .in1(R9702));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9884 (.out1(R9885), .clock(clock), .in1(R9884));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10011 (.out1(R10012), .clock(clock), .in1(R10011));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10133 (.out1(R10134), .clock(clock), .in1(R10133));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10302 (.out1(R10303), .clock(clock), .in1(R10302));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10415 (.out1(R10416), .clock(clock), .in1(R10415));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10523 (.out1(R10524), .clock(clock), .in1(R10523));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10679 (.out1(R10680), .clock(clock), .in1(R10679));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10779 (.out1(R10780), .clock(clock), .in1(R10779));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10874 (.out1(R10875), .clock(clock), .in1(R10874));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11016 (.out1(R11017), .clock(clock), .in1(R11016));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11103 (.out1(R11104), .clock(clock), .in1(_1155));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op1188 (.out1(_1150), .in1(ip2_3602_D), .in2(6 'd 34));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1189 (.out1(_1151), .in1(_1150));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op1190 (.out1(off_3635), .in1(_1151), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1195 (.out1(_1156), .in1(R11104), .in2(off_3635));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3850 (.out1(R3851), .clock(clock), .in1(R3850));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4106 (.out1(R4107), .clock(clock), .in1(R4106));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4361 (.out1(R4362), .clock(clock), .in1(R4361));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4606 (.out1(R4607), .clock(clock), .in1(R4606));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4846 (.out1(R4847), .clock(clock), .in1(R4846));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5133 (.out1(R5134), .clock(clock), .in1(R5133));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5365 (.out1(R5366), .clock(clock), .in1(R5365));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5592 (.out1(R5593), .clock(clock), .in1(R5592));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5866 (.out1(R5867), .clock(clock), .in1(R5866));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6084 (.out1(R6085), .clock(clock), .in1(R6084));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6297 (.out1(R6298), .clock(clock), .in1(R6297));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6558 (.out1(R6559), .clock(clock), .in1(R6558));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6763 (.out1(R6764), .clock(clock), .in1(R6763));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6963 (.out1(R6964), .clock(clock), .in1(R6963));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7210 (.out1(R7211), .clock(clock), .in1(R7210));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7402 (.out1(R7403), .clock(clock), .in1(R7402));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7589 (.out1(R7590), .clock(clock), .in1(R7589));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7823 (.out1(R7824), .clock(clock), .in1(R7823));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8002 (.out1(R8003), .clock(clock), .in1(R8002));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8176 (.out1(R8177), .clock(clock), .in1(R8176));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8397 (.out1(R8398), .clock(clock), .in1(R8397));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8563 (.out1(R8564), .clock(clock), .in1(R8563));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8724 (.out1(R8725), .clock(clock), .in1(R8724));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8932 (.out1(R8933), .clock(clock), .in1(R8932));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9085 (.out1(R9086), .clock(clock), .in1(R9085));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9233 (.out1(R9234), .clock(clock), .in1(R9233));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9428 (.out1(R9429), .clock(clock), .in1(R9428));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9568 (.out1(R9569), .clock(clock), .in1(R9568));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9703 (.out1(R9704), .clock(clock), .in1(R9703));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9885 (.out1(R9886), .clock(clock), .in1(R9885));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10012 (.out1(R10013), .clock(clock), .in1(R10012));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10134 (.out1(R10135), .clock(clock), .in1(R10134));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10303 (.out1(R10304), .clock(clock), .in1(R10303));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10416 (.out1(R10417), .clock(clock), .in1(R10416));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10524 (.out1(R10525), .clock(clock), .in1(R10524));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10680 (.out1(R10681), .clock(clock), .in1(R10680));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10780 (.out1(R10781), .clock(clock), .in1(R10780));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10875 (.out1(R10876), .clock(clock), .in1(R10875));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11017 (.out1(R11018), .clock(clock), .in1(R11017));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11104 (.out1(R11105), .clock(clock), .in1(off_3635));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11186 (.out1(R11187), .clock(clock), .in1(_1156));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op1196 (.out1(_1157), .in1(R11187), .in2(1 'd 1));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op1197 (.out1(ifout1197), .in1(_1157), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1265 (.out1(_1225), .in1(R11018));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1258 (.out1(_1218), .in1(R11018));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1247 (.out1(_1207), .in1(R11018));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1227 (.out1(_1187), .in1(R11018));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1266 (.out1(_1226), .in1(_1225), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1259 (.out1(_1219), .in1(_1218), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1248 (.out1(_1208), .in1(_1207), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1228 (.out1(_1188), .in1(_1187), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3851 (.out1(R3852), .clock(clock), .in1(R3851));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4107 (.out1(R4108), .clock(clock), .in1(R4107));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4362 (.out1(R4363), .clock(clock), .in1(R4362));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4607 (.out1(R4608), .clock(clock), .in1(R4607));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4847 (.out1(R4848), .clock(clock), .in1(R4847));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5134 (.out1(R5135), .clock(clock), .in1(R5134));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5366 (.out1(R5367), .clock(clock), .in1(R5366));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5593 (.out1(R5594), .clock(clock), .in1(R5593));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5867 (.out1(R5868), .clock(clock), .in1(R5867));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6085 (.out1(R6086), .clock(clock), .in1(R6085));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6298 (.out1(R6299), .clock(clock), .in1(R6298));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6559 (.out1(R6560), .clock(clock), .in1(R6559));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6764 (.out1(R6765), .clock(clock), .in1(R6764));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6964 (.out1(R6965), .clock(clock), .in1(R6964));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7211 (.out1(R7212), .clock(clock), .in1(R7211));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7403 (.out1(R7404), .clock(clock), .in1(R7403));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7590 (.out1(R7591), .clock(clock), .in1(R7590));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7824 (.out1(R7825), .clock(clock), .in1(R7824));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8003 (.out1(R8004), .clock(clock), .in1(R8003));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8177 (.out1(R8178), .clock(clock), .in1(R8177));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8398 (.out1(R8399), .clock(clock), .in1(R8398));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8564 (.out1(R8565), .clock(clock), .in1(R8564));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8725 (.out1(R8726), .clock(clock), .in1(R8725));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8933 (.out1(R8934), .clock(clock), .in1(R8933));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9086 (.out1(R9087), .clock(clock), .in1(R9086));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9234 (.out1(R9235), .clock(clock), .in1(R9234));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9429 (.out1(R9430), .clock(clock), .in1(R9429));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9569 (.out1(R9570), .clock(clock), .in1(R9569));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9704 (.out1(R9705), .clock(clock), .in1(R9704));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9886 (.out1(R9887), .clock(clock), .in1(R9886));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10013 (.out1(R10014), .clock(clock), .in1(R10013));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10135 (.out1(R10136), .clock(clock), .in1(R10135));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10304 (.out1(R10305), .clock(clock), .in1(R10304));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10417 (.out1(R10418), .clock(clock), .in1(R10417));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10525 (.out1(R10526), .clock(clock), .in1(R10525));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10681 (.out1(R10682), .clock(clock), .in1(R10681));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10781 (.out1(R10782), .clock(clock), .in1(R10781));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10876 (.out1(R10877), .clock(clock), .in1(R10876));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11018 (.out1(R11019), .clock(clock), .in1(R11018));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11105 (.out1(R11106), .clock(clock), .in1(R11105));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11187 (.out1(R11188), .clock(clock), .in1(ifout1197));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11276 (.out1(R11277), .clock(clock), .in1(_1226));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11277 (.out1(R11278), .clock(clock), .in1(_1219));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11278 (.out1(R11279), .clock(clock), .in1(_1208));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11279 (.out1(R11280), .clock(clock), .in1(_1188));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1240 (.out1(_1200), .in1(R11019));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1220 (.out1(_1180), .in1(R11019));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1209 (.out1(_1169), .in1(R11019));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1202 (.out1(_1162), .in1(R11019));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1269 (.out1(_1229), .in1(2 'd 2), .in2(R11106));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1241 (.out1(_1201), .in1(_1200), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1221 (.out1(_1181), .in1(_1180), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1210 (.out1(_1170), .in1(_1169), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1203 (.out1(_1163), .in1(_1162), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1267 (.out1(_1227), .in1(vec88_3636_D), .in2(R11277));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1260 (.out1(_1220), .in1(vec88_3636_D), .in2(R11278));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1249 (.out1(_1209), .in1(vec88_3636_D), .in2(R11279));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1229 (.out1(_1189), .in1(vec88_3636_D), .in2(R11280));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3852 (.out1(R3853), .clock(clock), .in1(R3852));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4108 (.out1(R4109), .clock(clock), .in1(R4108));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4363 (.out1(R4364), .clock(clock), .in1(R4363));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4608 (.out1(R4609), .clock(clock), .in1(R4608));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4848 (.out1(R4849), .clock(clock), .in1(R4848));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5135 (.out1(R5136), .clock(clock), .in1(R5135));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5367 (.out1(R5368), .clock(clock), .in1(R5367));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5594 (.out1(R5595), .clock(clock), .in1(R5594));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5868 (.out1(R5869), .clock(clock), .in1(R5868));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6086 (.out1(R6087), .clock(clock), .in1(R6086));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6299 (.out1(R6300), .clock(clock), .in1(R6299));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6560 (.out1(R6561), .clock(clock), .in1(R6560));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6765 (.out1(R6766), .clock(clock), .in1(R6765));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6965 (.out1(R6966), .clock(clock), .in1(R6965));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7212 (.out1(R7213), .clock(clock), .in1(R7212));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7404 (.out1(R7405), .clock(clock), .in1(R7404));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7591 (.out1(R7592), .clock(clock), .in1(R7591));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7825 (.out1(R7826), .clock(clock), .in1(R7825));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8004 (.out1(R8005), .clock(clock), .in1(R8004));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8178 (.out1(R8179), .clock(clock), .in1(R8178));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8399 (.out1(R8400), .clock(clock), .in1(R8399));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8565 (.out1(R8566), .clock(clock), .in1(R8565));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8726 (.out1(R8727), .clock(clock), .in1(R8726));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8934 (.out1(R8935), .clock(clock), .in1(R8934));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9087 (.out1(R9088), .clock(clock), .in1(R9087));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9235 (.out1(R9236), .clock(clock), .in1(R9235));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9430 (.out1(R9431), .clock(clock), .in1(R9430));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9570 (.out1(R9571), .clock(clock), .in1(R9570));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9705 (.out1(R9706), .clock(clock), .in1(R9705));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9887 (.out1(R9888), .clock(clock), .in1(R9887));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10014 (.out1(R10015), .clock(clock), .in1(R10014));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10136 (.out1(R10137), .clock(clock), .in1(R10136));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10305 (.out1(R10306), .clock(clock), .in1(R10305));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10418 (.out1(R10419), .clock(clock), .in1(R10418));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10526 (.out1(R10527), .clock(clock), .in1(R10526));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10682 (.out1(R10683), .clock(clock), .in1(R10682));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10782 (.out1(R10783), .clock(clock), .in1(R10782));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10877 (.out1(R10878), .clock(clock), .in1(R10877));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11019 (.out1(R11020), .clock(clock), .in1(R11019));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11106 (.out1(R11107), .clock(clock), .in1(R11106));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11188 (.out1(R11189), .clock(clock), .in1(R11188));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11280 (.out1(R11281), .clock(clock), .in1(_1229));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11281 (.out1(R11282), .clock(clock), .in1(_1201));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11282 (.out1(R11283), .clock(clock), .in1(_1181));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11283 (.out1(R11284), .clock(clock), .in1(_1170));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11284 (.out1(R11285), .clock(clock), .in1(_1163));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11285 (.out1(R11286), .clock(clock), .in1(_1227));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11286 (.out1(R11287), .clock(clock), .in1(_1220));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11287 (.out1(R11288), .clock(clock), .in1(_1209));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11288 (.out1(R11289), .clock(clock), .in1(_1189));
  SRAM op1268 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1228),.ADR(R11286));
  SRAM op1261 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1221),.ADR(R11287));
  SRAM op1250 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1210),.ADR(R11288));
  SRAM op1230 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1190),.ADR(R11289));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1262 (.out1(_1222), .in1(2 'd 2), .in2(R11107));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1251 (.out1(_1211), .in1(2 'd 2), .in2(R11107));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1244 (.out1(_1204), .in1(2 'd 2), .in2(R11107));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1231 (.out1(_1191), .in1(2 'd 2), .in2(R11107));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1224 (.out1(_1184), .in1(2 'd 2), .in2(R11107));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1213 (.out1(_1173), .in1(2 'd 2), .in2(R11107));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1242 (.out1(_1202), .in1(vec88_3636_D), .in2(R11282));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1222 (.out1(_1182), .in1(vec88_3636_D), .in2(R11283));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1211 (.out1(_1171), .in1(vec88_3636_D), .in2(R11284));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1204 (.out1(_1164), .in1(vec88_3636_D), .in2(R11285));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1270 (.out1(_1230), .in1(R11281), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3853 (.out1(R3854), .clock(clock), .in1(R3853));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4109 (.out1(R4110), .clock(clock), .in1(R4109));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4364 (.out1(R4365), .clock(clock), .in1(R4364));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4609 (.out1(R4610), .clock(clock), .in1(R4609));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4849 (.out1(R4850), .clock(clock), .in1(R4849));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5136 (.out1(R5137), .clock(clock), .in1(R5136));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5368 (.out1(R5369), .clock(clock), .in1(R5368));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5595 (.out1(R5596), .clock(clock), .in1(R5595));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5869 (.out1(R5870), .clock(clock), .in1(R5869));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6087 (.out1(R6088), .clock(clock), .in1(R6087));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6300 (.out1(R6301), .clock(clock), .in1(R6300));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6561 (.out1(R6562), .clock(clock), .in1(R6561));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6766 (.out1(R6767), .clock(clock), .in1(R6766));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6966 (.out1(R6967), .clock(clock), .in1(R6966));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7213 (.out1(R7214), .clock(clock), .in1(R7213));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7405 (.out1(R7406), .clock(clock), .in1(R7405));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7592 (.out1(R7593), .clock(clock), .in1(R7592));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7826 (.out1(R7827), .clock(clock), .in1(R7826));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8005 (.out1(R8006), .clock(clock), .in1(R8005));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8179 (.out1(R8180), .clock(clock), .in1(R8179));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8400 (.out1(R8401), .clock(clock), .in1(R8400));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8566 (.out1(R8567), .clock(clock), .in1(R8566));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8727 (.out1(R8728), .clock(clock), .in1(R8727));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8935 (.out1(R8936), .clock(clock), .in1(R8935));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9088 (.out1(R9089), .clock(clock), .in1(R9088));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9236 (.out1(R9237), .clock(clock), .in1(R9236));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9431 (.out1(R9432), .clock(clock), .in1(R9431));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9571 (.out1(R9572), .clock(clock), .in1(R9571));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9706 (.out1(R9707), .clock(clock), .in1(R9706));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9888 (.out1(R9889), .clock(clock), .in1(R9888));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10015 (.out1(R10016), .clock(clock), .in1(R10015));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10137 (.out1(R10138), .clock(clock), .in1(R10137));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10306 (.out1(R10307), .clock(clock), .in1(R10306));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10419 (.out1(R10420), .clock(clock), .in1(R10419));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10527 (.out1(R10528), .clock(clock), .in1(R10527));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10683 (.out1(R10684), .clock(clock), .in1(R10683));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10783 (.out1(R10784), .clock(clock), .in1(R10783));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10878 (.out1(R10879), .clock(clock), .in1(R10878));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11020 (.out1(R11021), .clock(clock), .in1(R11020));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11107 (.out1(R11108), .clock(clock), .in1(R11107));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11189 (.out1(R11190), .clock(clock), .in1(R11189));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11289 (.out1(R11290), .clock(clock), .in1(_1228));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11290 (.out1(R11291), .clock(clock), .in1(_1221));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11291 (.out1(R11292), .clock(clock), .in1(_1210));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11292 (.out1(R11293), .clock(clock), .in1(_1190));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11293 (.out1(R11294), .clock(clock), .in1(_1222));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11294 (.out1(R11295), .clock(clock), .in1(_1211));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11295 (.out1(R11296), .clock(clock), .in1(_1204));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11296 (.out1(R11297), .clock(clock), .in1(_1191));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11297 (.out1(R11298), .clock(clock), .in1(_1184));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11298 (.out1(R11299), .clock(clock), .in1(_1173));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11299 (.out1(R11300), .clock(clock), .in1(_1202));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11300 (.out1(R11301), .clock(clock), .in1(_1182));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11301 (.out1(R11302), .clock(clock), .in1(_1171));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11302 (.out1(R11303), .clock(clock), .in1(_1164));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11303 (.out1(R11304), .clock(clock), .in1(_1230));
  SRAM op1243 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1203),.ADR(R11300));
  SRAM op1223 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1183),.ADR(R11301));
  SRAM op1212 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1172),.ADR(R11302));
  SRAM op1205 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1165),.ADR(R11303));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1271 (.out1(_1231), .in1(R11290), .in2(R11304));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1272 (.out1(_1232), .in1(_1231), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1263 (.out1(_1223), .in1(R11294), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1252 (.out1(_1212), .in1(R11295), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1232 (.out1(_1192), .in1(R11297), .in2(64 'd 18446744073709551615));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1206 (.out1(_1166), .in1(2 'd 2), .in2(R11108));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1273 (.out1(_1233), .in1(_1232), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1264 (.out1(_1224), .in1(R11291), .in2(_1223));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1253 (.out1(_1213), .in1(R11292), .in2(_1212));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1233 (.out1(_1193), .in1(R11293), .in2(_1192));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1274 (.out1(_1234), .in1(_1224), .in2(_1233));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1254 (.out1(_1214), .in1(_1213), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1245 (.out1(_1205), .in1(R11296), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1234 (.out1(_1194), .in1(_1193), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1225 (.out1(_1185), .in1(R11298), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1214 (.out1(_1174), .in1(R11299), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3854 (.out1(R3855), .clock(clock), .in1(R3854));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4110 (.out1(R4111), .clock(clock), .in1(R4110));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4365 (.out1(R4366), .clock(clock), .in1(R4365));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4610 (.out1(R4611), .clock(clock), .in1(R4610));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4850 (.out1(R4851), .clock(clock), .in1(R4850));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5137 (.out1(R5138), .clock(clock), .in1(R5137));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5369 (.out1(R5370), .clock(clock), .in1(R5369));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5596 (.out1(R5597), .clock(clock), .in1(R5596));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5870 (.out1(R5871), .clock(clock), .in1(R5870));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6088 (.out1(R6089), .clock(clock), .in1(R6088));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6301 (.out1(R6302), .clock(clock), .in1(R6301));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6562 (.out1(R6563), .clock(clock), .in1(R6562));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6767 (.out1(R6768), .clock(clock), .in1(R6767));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6967 (.out1(R6968), .clock(clock), .in1(R6967));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7214 (.out1(R7215), .clock(clock), .in1(R7214));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7406 (.out1(R7407), .clock(clock), .in1(R7406));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7593 (.out1(R7594), .clock(clock), .in1(R7593));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7827 (.out1(R7828), .clock(clock), .in1(R7827));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8006 (.out1(R8007), .clock(clock), .in1(R8006));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8180 (.out1(R8181), .clock(clock), .in1(R8180));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8401 (.out1(R8402), .clock(clock), .in1(R8401));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8567 (.out1(R8568), .clock(clock), .in1(R8567));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8728 (.out1(R8729), .clock(clock), .in1(R8728));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8936 (.out1(R8937), .clock(clock), .in1(R8936));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9089 (.out1(R9090), .clock(clock), .in1(R9089));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9237 (.out1(R9238), .clock(clock), .in1(R9237));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9432 (.out1(R9433), .clock(clock), .in1(R9432));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9572 (.out1(R9573), .clock(clock), .in1(R9572));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9707 (.out1(R9708), .clock(clock), .in1(R9707));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9889 (.out1(R9890), .clock(clock), .in1(R9889));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10016 (.out1(R10017), .clock(clock), .in1(R10016));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10138 (.out1(R10139), .clock(clock), .in1(R10138));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10307 (.out1(R10308), .clock(clock), .in1(R10307));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10420 (.out1(R10421), .clock(clock), .in1(R10420));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10528 (.out1(R10529), .clock(clock), .in1(R10528));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10684 (.out1(R10685), .clock(clock), .in1(R10684));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10784 (.out1(R10785), .clock(clock), .in1(R10784));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10879 (.out1(R10880), .clock(clock), .in1(R10879));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11021 (.out1(R11022), .clock(clock), .in1(R11021));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11108 (.out1(R11109), .clock(clock), .in1(R11108));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11190 (.out1(R11191), .clock(clock), .in1(R11190));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11304 (.out1(R11305), .clock(clock), .in1(_1203));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11305 (.out1(R11306), .clock(clock), .in1(_1183));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11306 (.out1(R11307), .clock(clock), .in1(_1172));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11307 (.out1(R11308), .clock(clock), .in1(_1165));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11308 (.out1(R11309), .clock(clock), .in1(_1166));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11309 (.out1(R11310), .clock(clock), .in1(_1234));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11310 (.out1(R11311), .clock(clock), .in1(_1214));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11311 (.out1(R11312), .clock(clock), .in1(_1205));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11312 (.out1(R11313), .clock(clock), .in1(_1194));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11313 (.out1(R11314), .clock(clock), .in1(_1185));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11314 (.out1(R11315), .clock(clock), .in1(_1174));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1255 (.out1(_1215), .in1(R11311), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1246 (.out1(_1206), .in1(R11305), .in2(R11312));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1215 (.out1(_1175), .in1(R11307), .in2(R11315));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1275 (.out1(_1235), .in1(R11310), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1256 (.out1(_1216), .in1(_1206), .in2(_1215));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1235 (.out1(_1195), .in1(R11313), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1226 (.out1(_1186), .in1(R11306), .in2(R11314));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1216 (.out1(_1176), .in1(_1175), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1207 (.out1(_1167), .in1(R11309), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1236 (.out1(_1196), .in1(_1186), .in2(_1195));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1276 (.out1(_1236), .in1(_1235), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1257 (.out1(_1217), .in1(_1216), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1217 (.out1(_1177), .in1(_1176), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1208 (.out1(_1168), .in1(R11308), .in2(_1167));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1277 (.out1(_1237), .in1(_1217), .in2(_1236));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1237 (.out1(_1197), .in1(_1196), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1218 (.out1(_1178), .in1(_1168), .in2(_1177));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3855 (.out1(R3856), .clock(clock), .in1(R3855));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4111 (.out1(R4112), .clock(clock), .in1(R4111));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4366 (.out1(R4367), .clock(clock), .in1(R4366));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4611 (.out1(R4612), .clock(clock), .in1(R4611));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4851 (.out1(R4852), .clock(clock), .in1(R4851));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5138 (.out1(R5139), .clock(clock), .in1(R5138));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5370 (.out1(R5371), .clock(clock), .in1(R5370));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5597 (.out1(R5598), .clock(clock), .in1(R5597));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5871 (.out1(R5872), .clock(clock), .in1(R5871));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6089 (.out1(R6090), .clock(clock), .in1(R6089));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6302 (.out1(R6303), .clock(clock), .in1(R6302));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6563 (.out1(R6564), .clock(clock), .in1(R6563));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6768 (.out1(R6769), .clock(clock), .in1(R6768));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6968 (.out1(R6969), .clock(clock), .in1(R6968));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7215 (.out1(R7216), .clock(clock), .in1(R7215));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7407 (.out1(R7408), .clock(clock), .in1(R7407));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7594 (.out1(R7595), .clock(clock), .in1(R7594));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7828 (.out1(R7829), .clock(clock), .in1(R7828));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8007 (.out1(R8008), .clock(clock), .in1(R8007));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8181 (.out1(R8182), .clock(clock), .in1(R8181));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8402 (.out1(R8403), .clock(clock), .in1(R8402));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8568 (.out1(R8569), .clock(clock), .in1(R8568));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8729 (.out1(R8730), .clock(clock), .in1(R8729));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8937 (.out1(R8938), .clock(clock), .in1(R8937));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9090 (.out1(R9091), .clock(clock), .in1(R9090));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9238 (.out1(R9239), .clock(clock), .in1(R9238));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9433 (.out1(R9434), .clock(clock), .in1(R9433));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9573 (.out1(R9574), .clock(clock), .in1(R9573));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9708 (.out1(R9709), .clock(clock), .in1(R9708));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9890 (.out1(R9891), .clock(clock), .in1(R9890));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10017 (.out1(R10018), .clock(clock), .in1(R10017));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10139 (.out1(R10140), .clock(clock), .in1(R10139));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10308 (.out1(R10309), .clock(clock), .in1(R10308));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10421 (.out1(R10422), .clock(clock), .in1(R10421));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10529 (.out1(R10530), .clock(clock), .in1(R10529));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10685 (.out1(R10686), .clock(clock), .in1(R10685));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10785 (.out1(R10786), .clock(clock), .in1(R10785));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10880 (.out1(R10881), .clock(clock), .in1(R10880));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11022 (.out1(R11023), .clock(clock), .in1(R11022));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11109 (.out1(R11110), .clock(clock), .in1(R11109));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11191 (.out1(R11192), .clock(clock), .in1(R11191));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11315 (.out1(R11316), .clock(clock), .in1(_1237));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11316 (.out1(R11317), .clock(clock), .in1(_1197));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11317 (.out1(R11318), .clock(clock), .in1(_1178));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1198 (.out1(_1158), .in1(R11023));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1238 (.out1(_1198), .in1(R11317), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1219 (.out1(_1179), .in1(R11318), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op1278 (.out1(_1238), .in1(R11316), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1239 (.out1(_1199), .in1(_1179), .in2(_1198));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1199 (.out1(_1159), .in1(_1158), .in2(2 'd 2));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1279 (.out1(_1239), .in1(_1199), .in2(_1238));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op1280 (.out1(_1240), .in1(_1239), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3856 (.out1(R3857), .clock(clock), .in1(R3856));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4112 (.out1(R4113), .clock(clock), .in1(R4112));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4367 (.out1(R4368), .clock(clock), .in1(R4367));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4612 (.out1(R4613), .clock(clock), .in1(R4612));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4852 (.out1(R4853), .clock(clock), .in1(R4852));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5139 (.out1(R5140), .clock(clock), .in1(R5139));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5371 (.out1(R5372), .clock(clock), .in1(R5371));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5598 (.out1(R5599), .clock(clock), .in1(R5598));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5872 (.out1(R5873), .clock(clock), .in1(R5872));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6090 (.out1(R6091), .clock(clock), .in1(R6090));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6303 (.out1(R6304), .clock(clock), .in1(R6303));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6564 (.out1(R6565), .clock(clock), .in1(R6564));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6769 (.out1(R6770), .clock(clock), .in1(R6769));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6969 (.out1(R6970), .clock(clock), .in1(R6969));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7216 (.out1(R7217), .clock(clock), .in1(R7216));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7408 (.out1(R7409), .clock(clock), .in1(R7408));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7595 (.out1(R7596), .clock(clock), .in1(R7595));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7829 (.out1(R7830), .clock(clock), .in1(R7829));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8008 (.out1(R8009), .clock(clock), .in1(R8008));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8182 (.out1(R8183), .clock(clock), .in1(R8182));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8403 (.out1(R8404), .clock(clock), .in1(R8403));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8569 (.out1(R8570), .clock(clock), .in1(R8569));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8730 (.out1(R8731), .clock(clock), .in1(R8730));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8938 (.out1(R8939), .clock(clock), .in1(R8938));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9091 (.out1(R9092), .clock(clock), .in1(R9091));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9239 (.out1(R9240), .clock(clock), .in1(R9239));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9434 (.out1(R9435), .clock(clock), .in1(R9434));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9574 (.out1(R9575), .clock(clock), .in1(R9574));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9709 (.out1(R9710), .clock(clock), .in1(R9709));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9891 (.out1(R9892), .clock(clock), .in1(R9891));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10018 (.out1(R10019), .clock(clock), .in1(R10018));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10140 (.out1(R10141), .clock(clock), .in1(R10140));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10309 (.out1(R10310), .clock(clock), .in1(R10309));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10422 (.out1(R10423), .clock(clock), .in1(R10422));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10530 (.out1(R10531), .clock(clock), .in1(R10530));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10686 (.out1(R10687), .clock(clock), .in1(R10686));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10786 (.out1(R10787), .clock(clock), .in1(R10786));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10881 (.out1(R10882), .clock(clock), .in1(R10881));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11023 (.out1(R11024), .clock(clock), .in1(R11023));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11110 (.out1(R11111), .clock(clock), .in1(R11110));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11192 (.out1(R11193), .clock(clock), .in1(R11192));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11318 (.out1(R11319), .clock(clock), .in1(_1159));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11319 (.out1(R11320), .clock(clock), .in1(_1240));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op1281 (.out1(_1241), .in1(R11320), .in2(57 'd 72340172838076673));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1200 (.out1(_1160), .in1(base0_88_3641_D), .in2(R11319));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3857 (.out1(R3858), .clock(clock), .in1(R3857));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4113 (.out1(R4114), .clock(clock), .in1(R4113));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4368 (.out1(R4369), .clock(clock), .in1(R4368));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4613 (.out1(R4614), .clock(clock), .in1(R4613));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4853 (.out1(R4854), .clock(clock), .in1(R4853));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5140 (.out1(R5141), .clock(clock), .in1(R5140));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5372 (.out1(R5373), .clock(clock), .in1(R5372));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5599 (.out1(R5600), .clock(clock), .in1(R5599));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5873 (.out1(R5874), .clock(clock), .in1(R5873));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6091 (.out1(R6092), .clock(clock), .in1(R6091));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6304 (.out1(R6305), .clock(clock), .in1(R6304));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6565 (.out1(R6566), .clock(clock), .in1(R6565));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6770 (.out1(R6771), .clock(clock), .in1(R6770));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6970 (.out1(R6971), .clock(clock), .in1(R6970));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7217 (.out1(R7218), .clock(clock), .in1(R7217));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7409 (.out1(R7410), .clock(clock), .in1(R7409));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7596 (.out1(R7597), .clock(clock), .in1(R7596));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7830 (.out1(R7831), .clock(clock), .in1(R7830));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8009 (.out1(R8010), .clock(clock), .in1(R8009));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8183 (.out1(R8184), .clock(clock), .in1(R8183));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8404 (.out1(R8405), .clock(clock), .in1(R8404));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8570 (.out1(R8571), .clock(clock), .in1(R8570));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8731 (.out1(R8732), .clock(clock), .in1(R8731));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8939 (.out1(R8940), .clock(clock), .in1(R8939));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9092 (.out1(R9093), .clock(clock), .in1(R9092));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9240 (.out1(R9241), .clock(clock), .in1(R9240));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9435 (.out1(R9436), .clock(clock), .in1(R9435));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9575 (.out1(R9576), .clock(clock), .in1(R9575));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9710 (.out1(R9711), .clock(clock), .in1(R9710));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9892 (.out1(R9893), .clock(clock), .in1(R9892));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10019 (.out1(R10020), .clock(clock), .in1(R10019));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10141 (.out1(R10142), .clock(clock), .in1(R10141));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10310 (.out1(R10311), .clock(clock), .in1(R10310));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10423 (.out1(R10424), .clock(clock), .in1(R10423));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10531 (.out1(R10532), .clock(clock), .in1(R10531));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10687 (.out1(R10688), .clock(clock), .in1(R10687));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10787 (.out1(R10788), .clock(clock), .in1(R10787));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10882 (.out1(R10883), .clock(clock), .in1(R10882));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11024 (.out1(R11025), .clock(clock), .in1(R11024));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11111 (.out1(R11112), .clock(clock), .in1(R11111));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11193 (.out1(R11194), .clock(clock), .in1(R11193));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11320 (.out1(R11321), .clock(clock), .in1(_1241));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11321 (.out1(R11322), .clock(clock), .in1(_1160));
  SRAM op1201 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1161),.ADR(R11322));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op1282 (.out1(_1242), .in1(R11321), .in2(6 'd 56));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3858 (.out1(R3859), .clock(clock), .in1(R3858));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4114 (.out1(R4115), .clock(clock), .in1(R4114));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4369 (.out1(R4370), .clock(clock), .in1(R4369));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4614 (.out1(R4615), .clock(clock), .in1(R4614));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4854 (.out1(R4855), .clock(clock), .in1(R4854));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5141 (.out1(R5142), .clock(clock), .in1(R5141));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5373 (.out1(R5374), .clock(clock), .in1(R5373));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5600 (.out1(R5601), .clock(clock), .in1(R5600));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5874 (.out1(R5875), .clock(clock), .in1(R5874));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6092 (.out1(R6093), .clock(clock), .in1(R6092));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6305 (.out1(R6306), .clock(clock), .in1(R6305));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6566 (.out1(R6567), .clock(clock), .in1(R6566));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6771 (.out1(R6772), .clock(clock), .in1(R6771));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6971 (.out1(R6972), .clock(clock), .in1(R6971));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7218 (.out1(R7219), .clock(clock), .in1(R7218));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7410 (.out1(R7411), .clock(clock), .in1(R7410));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7597 (.out1(R7598), .clock(clock), .in1(R7597));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7831 (.out1(R7832), .clock(clock), .in1(R7831));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8010 (.out1(R8011), .clock(clock), .in1(R8010));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8184 (.out1(R8185), .clock(clock), .in1(R8184));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8405 (.out1(R8406), .clock(clock), .in1(R8405));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8571 (.out1(R8572), .clock(clock), .in1(R8571));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8732 (.out1(R8733), .clock(clock), .in1(R8732));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8940 (.out1(R8941), .clock(clock), .in1(R8940));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9093 (.out1(R9094), .clock(clock), .in1(R9093));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9241 (.out1(R9242), .clock(clock), .in1(R9241));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9436 (.out1(R9437), .clock(clock), .in1(R9436));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9576 (.out1(R9577), .clock(clock), .in1(R9576));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9711 (.out1(R9712), .clock(clock), .in1(R9711));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9893 (.out1(R9894), .clock(clock), .in1(R9893));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10020 (.out1(R10021), .clock(clock), .in1(R10020));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10142 (.out1(R10143), .clock(clock), .in1(R10142));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10311 (.out1(R10312), .clock(clock), .in1(R10311));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10424 (.out1(R10425), .clock(clock), .in1(R10424));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10532 (.out1(R10533), .clock(clock), .in1(R10532));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10688 (.out1(R10689), .clock(clock), .in1(R10688));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10788 (.out1(R10789), .clock(clock), .in1(R10788));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10883 (.out1(R10884), .clock(clock), .in1(R10883));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11025 (.out1(R11026), .clock(clock), .in1(R11025));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11112 (.out1(R11113), .clock(clock), .in1(R11112));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11194 (.out1(R11195), .clock(clock), .in1(R11194));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11322 (.out1(R11323), .clock(clock), .in1(_1161));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11323 (.out1(R11324), .clock(clock), .in1(_1242));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1283 (.out1(_1243), .in1(R11324));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1284 (.out1(_1244), .in1(R11323), .in2(_1243));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1285 (.out1(idx_3642), .in1(_1244), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3859 (.out1(R3860), .clock(clock), .in1(R3859));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4115 (.out1(R4116), .clock(clock), .in1(R4115));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4370 (.out1(R4371), .clock(clock), .in1(R4370));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4615 (.out1(R4616), .clock(clock), .in1(R4615));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4855 (.out1(R4856), .clock(clock), .in1(R4855));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5142 (.out1(R5143), .clock(clock), .in1(R5142));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5374 (.out1(R5375), .clock(clock), .in1(R5374));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5601 (.out1(R5602), .clock(clock), .in1(R5601));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5875 (.out1(R5876), .clock(clock), .in1(R5875));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6093 (.out1(R6094), .clock(clock), .in1(R6093));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6306 (.out1(R6307), .clock(clock), .in1(R6306));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6567 (.out1(R6568), .clock(clock), .in1(R6567));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6772 (.out1(R6773), .clock(clock), .in1(R6772));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6972 (.out1(R6973), .clock(clock), .in1(R6972));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7219 (.out1(R7220), .clock(clock), .in1(R7219));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7411 (.out1(R7412), .clock(clock), .in1(R7411));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7598 (.out1(R7599), .clock(clock), .in1(R7598));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7832 (.out1(R7833), .clock(clock), .in1(R7832));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8011 (.out1(R8012), .clock(clock), .in1(R8011));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8185 (.out1(R8186), .clock(clock), .in1(R8185));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8406 (.out1(R8407), .clock(clock), .in1(R8406));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8572 (.out1(R8573), .clock(clock), .in1(R8572));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8733 (.out1(R8734), .clock(clock), .in1(R8733));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8941 (.out1(R8942), .clock(clock), .in1(R8941));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9094 (.out1(R9095), .clock(clock), .in1(R9094));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9242 (.out1(R9243), .clock(clock), .in1(R9242));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9437 (.out1(R9438), .clock(clock), .in1(R9437));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9577 (.out1(R9578), .clock(clock), .in1(R9577));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9712 (.out1(R9713), .clock(clock), .in1(R9712));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9894 (.out1(R9895), .clock(clock), .in1(R9894));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10021 (.out1(R10022), .clock(clock), .in1(R10021));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10143 (.out1(R10144), .clock(clock), .in1(R10143));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10312 (.out1(R10313), .clock(clock), .in1(R10312));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10425 (.out1(R10426), .clock(clock), .in1(R10425));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10533 (.out1(R10534), .clock(clock), .in1(R10533));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10689 (.out1(R10690), .clock(clock), .in1(R10689));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10789 (.out1(R10790), .clock(clock), .in1(R10789));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10884 (.out1(R10885), .clock(clock), .in1(R10884));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11026 (.out1(R11027), .clock(clock), .in1(R11026));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11113 (.out1(R11114), .clock(clock), .in1(R11113));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11195 (.out1(R11196), .clock(clock), .in1(R11195));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11324 (.out1(R11325), .clock(clock), .in1(idx_3642));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1289 (.out1(_1247), .in1(R11325));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1290 (.out1(_1248), .in1(_1247), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3860 (.out1(R3861), .clock(clock), .in1(R3860));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4116 (.out1(R4117), .clock(clock), .in1(R4116));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4371 (.out1(R4372), .clock(clock), .in1(R4371));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4616 (.out1(R4617), .clock(clock), .in1(R4616));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4856 (.out1(R4857), .clock(clock), .in1(R4856));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5143 (.out1(R5144), .clock(clock), .in1(R5143));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5375 (.out1(R5376), .clock(clock), .in1(R5375));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5602 (.out1(R5603), .clock(clock), .in1(R5602));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5876 (.out1(R5877), .clock(clock), .in1(R5876));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6094 (.out1(R6095), .clock(clock), .in1(R6094));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6307 (.out1(R6308), .clock(clock), .in1(R6307));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6568 (.out1(R6569), .clock(clock), .in1(R6568));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6773 (.out1(R6774), .clock(clock), .in1(R6773));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6973 (.out1(R6974), .clock(clock), .in1(R6973));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7220 (.out1(R7221), .clock(clock), .in1(R7220));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7412 (.out1(R7413), .clock(clock), .in1(R7412));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7599 (.out1(R7600), .clock(clock), .in1(R7599));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7833 (.out1(R7834), .clock(clock), .in1(R7833));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8012 (.out1(R8013), .clock(clock), .in1(R8012));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8186 (.out1(R8187), .clock(clock), .in1(R8186));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8407 (.out1(R8408), .clock(clock), .in1(R8407));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8573 (.out1(R8574), .clock(clock), .in1(R8573));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8734 (.out1(R8735), .clock(clock), .in1(R8734));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8942 (.out1(R8943), .clock(clock), .in1(R8942));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9095 (.out1(R9096), .clock(clock), .in1(R9095));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9243 (.out1(R9244), .clock(clock), .in1(R9243));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9438 (.out1(R9439), .clock(clock), .in1(R9438));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9578 (.out1(R9579), .clock(clock), .in1(R9578));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9713 (.out1(R9714), .clock(clock), .in1(R9713));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9895 (.out1(R9896), .clock(clock), .in1(R9895));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10022 (.out1(R10023), .clock(clock), .in1(R10022));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10144 (.out1(R10145), .clock(clock), .in1(R10144));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10313 (.out1(R10314), .clock(clock), .in1(R10313));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10426 (.out1(R10427), .clock(clock), .in1(R10426));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10534 (.out1(R10535), .clock(clock), .in1(R10534));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10690 (.out1(R10691), .clock(clock), .in1(R10690));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10790 (.out1(R10791), .clock(clock), .in1(R10790));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10885 (.out1(R10886), .clock(clock), .in1(R10885));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11027 (.out1(R11028), .clock(clock), .in1(R11027));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11114 (.out1(R11115), .clock(clock), .in1(R11114));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11196 (.out1(R11197), .clock(clock), .in1(R11196));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11325 (.out1(R11326), .clock(clock), .in1(R11325));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11399 (.out1(R11400), .clock(clock), .in1(_1248));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1291 (.out1(_1249), .in1(vec94_3644_D), .in2(R11400));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3861 (.out1(R3862), .clock(clock), .in1(R3861));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4117 (.out1(R4118), .clock(clock), .in1(R4117));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4372 (.out1(R4373), .clock(clock), .in1(R4372));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4617 (.out1(R4618), .clock(clock), .in1(R4617));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4857 (.out1(R4858), .clock(clock), .in1(R4857));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5144 (.out1(R5145), .clock(clock), .in1(R5144));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5376 (.out1(R5377), .clock(clock), .in1(R5376));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5603 (.out1(R5604), .clock(clock), .in1(R5603));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5877 (.out1(R5878), .clock(clock), .in1(R5877));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6095 (.out1(R6096), .clock(clock), .in1(R6095));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6308 (.out1(R6309), .clock(clock), .in1(R6308));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6569 (.out1(R6570), .clock(clock), .in1(R6569));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6774 (.out1(R6775), .clock(clock), .in1(R6774));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6974 (.out1(R6975), .clock(clock), .in1(R6974));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7221 (.out1(R7222), .clock(clock), .in1(R7221));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7413 (.out1(R7414), .clock(clock), .in1(R7413));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7600 (.out1(R7601), .clock(clock), .in1(R7600));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7834 (.out1(R7835), .clock(clock), .in1(R7834));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8013 (.out1(R8014), .clock(clock), .in1(R8013));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8187 (.out1(R8188), .clock(clock), .in1(R8187));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8408 (.out1(R8409), .clock(clock), .in1(R8408));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8574 (.out1(R8575), .clock(clock), .in1(R8574));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8735 (.out1(R8736), .clock(clock), .in1(R8735));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8943 (.out1(R8944), .clock(clock), .in1(R8943));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9096 (.out1(R9097), .clock(clock), .in1(R9096));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9244 (.out1(R9245), .clock(clock), .in1(R9244));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9439 (.out1(R9440), .clock(clock), .in1(R9439));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9579 (.out1(R9580), .clock(clock), .in1(R9579));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9714 (.out1(R9715), .clock(clock), .in1(R9714));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9896 (.out1(R9897), .clock(clock), .in1(R9896));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10023 (.out1(R10024), .clock(clock), .in1(R10023));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10145 (.out1(R10146), .clock(clock), .in1(R10145));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10314 (.out1(R10315), .clock(clock), .in1(R10314));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10427 (.out1(R10428), .clock(clock), .in1(R10427));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10535 (.out1(R10536), .clock(clock), .in1(R10535));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10691 (.out1(R10692), .clock(clock), .in1(R10691));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10791 (.out1(R10792), .clock(clock), .in1(R10791));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10886 (.out1(R10887), .clock(clock), .in1(R10886));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11028 (.out1(R11029), .clock(clock), .in1(R11028));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11115 (.out1(R11116), .clock(clock), .in1(R11115));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11197 (.out1(R11198), .clock(clock), .in1(R11197));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11326 (.out1(R11327), .clock(clock), .in1(R11326));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11400 (.out1(R11401), .clock(clock), .in1(_1249));
  SRAM op1292 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1250),.ADR(R11401));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3862 (.out1(R3863), .clock(clock), .in1(R3862));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4118 (.out1(R4119), .clock(clock), .in1(R4118));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4373 (.out1(R4374), .clock(clock), .in1(R4373));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4618 (.out1(R4619), .clock(clock), .in1(R4618));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4858 (.out1(R4859), .clock(clock), .in1(R4858));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5145 (.out1(R5146), .clock(clock), .in1(R5145));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5377 (.out1(R5378), .clock(clock), .in1(R5377));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5604 (.out1(R5605), .clock(clock), .in1(R5604));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5878 (.out1(R5879), .clock(clock), .in1(R5878));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6096 (.out1(R6097), .clock(clock), .in1(R6096));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6309 (.out1(R6310), .clock(clock), .in1(R6309));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6570 (.out1(R6571), .clock(clock), .in1(R6570));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6775 (.out1(R6776), .clock(clock), .in1(R6775));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6975 (.out1(R6976), .clock(clock), .in1(R6975));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7222 (.out1(R7223), .clock(clock), .in1(R7222));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7414 (.out1(R7415), .clock(clock), .in1(R7414));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7601 (.out1(R7602), .clock(clock), .in1(R7601));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7835 (.out1(R7836), .clock(clock), .in1(R7835));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8014 (.out1(R8015), .clock(clock), .in1(R8014));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8188 (.out1(R8189), .clock(clock), .in1(R8188));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8409 (.out1(R8410), .clock(clock), .in1(R8409));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8575 (.out1(R8576), .clock(clock), .in1(R8575));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8736 (.out1(R8737), .clock(clock), .in1(R8736));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8944 (.out1(R8945), .clock(clock), .in1(R8944));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9097 (.out1(R9098), .clock(clock), .in1(R9097));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9245 (.out1(R9246), .clock(clock), .in1(R9245));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9440 (.out1(R9441), .clock(clock), .in1(R9440));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9580 (.out1(R9581), .clock(clock), .in1(R9580));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9715 (.out1(R9716), .clock(clock), .in1(R9715));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9897 (.out1(R9898), .clock(clock), .in1(R9897));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10024 (.out1(R10025), .clock(clock), .in1(R10024));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10146 (.out1(R10147), .clock(clock), .in1(R10146));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10315 (.out1(R10316), .clock(clock), .in1(R10315));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10428 (.out1(R10429), .clock(clock), .in1(R10428));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10536 (.out1(R10537), .clock(clock), .in1(R10536));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10692 (.out1(R10693), .clock(clock), .in1(R10692));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10792 (.out1(R10793), .clock(clock), .in1(R10792));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10887 (.out1(R10888), .clock(clock), .in1(R10887));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11029 (.out1(R11030), .clock(clock), .in1(R11029));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11116 (.out1(R11117), .clock(clock), .in1(R11116));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11198 (.out1(R11199), .clock(clock), .in1(R11198));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11327 (.out1(R11328), .clock(clock), .in1(R11327));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11401 (.out1(R11402), .clock(clock), .in1(_1250));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(5), .BITSIZE_out1(64), .PRECISION(64)) op1286 (.out1(_1245), .in1(ip2_3602_D), .in2(5 'd 28));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1287 (.out1(_1246), .in1(_1245));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op1288 (.out1(off_3643), .in1(_1246), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1293 (.out1(_1251), .in1(R11402), .in2(off_3643));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3863 (.out1(R3864), .clock(clock), .in1(R3863));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4119 (.out1(R4120), .clock(clock), .in1(R4119));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4374 (.out1(R4375), .clock(clock), .in1(R4374));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4619 (.out1(R4620), .clock(clock), .in1(R4619));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4859 (.out1(R4860), .clock(clock), .in1(R4859));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5146 (.out1(R5147), .clock(clock), .in1(R5146));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5378 (.out1(R5379), .clock(clock), .in1(R5378));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5605 (.out1(R5606), .clock(clock), .in1(R5605));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5879 (.out1(R5880), .clock(clock), .in1(R5879));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6097 (.out1(R6098), .clock(clock), .in1(R6097));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6310 (.out1(R6311), .clock(clock), .in1(R6310));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6571 (.out1(R6572), .clock(clock), .in1(R6571));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6776 (.out1(R6777), .clock(clock), .in1(R6776));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6976 (.out1(R6977), .clock(clock), .in1(R6976));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7223 (.out1(R7224), .clock(clock), .in1(R7223));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7415 (.out1(R7416), .clock(clock), .in1(R7415));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7602 (.out1(R7603), .clock(clock), .in1(R7602));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7836 (.out1(R7837), .clock(clock), .in1(R7836));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8015 (.out1(R8016), .clock(clock), .in1(R8015));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8189 (.out1(R8190), .clock(clock), .in1(R8189));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8410 (.out1(R8411), .clock(clock), .in1(R8410));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8576 (.out1(R8577), .clock(clock), .in1(R8576));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8737 (.out1(R8738), .clock(clock), .in1(R8737));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8945 (.out1(R8946), .clock(clock), .in1(R8945));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9098 (.out1(R9099), .clock(clock), .in1(R9098));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9246 (.out1(R9247), .clock(clock), .in1(R9246));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9441 (.out1(R9442), .clock(clock), .in1(R9441));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9581 (.out1(R9582), .clock(clock), .in1(R9581));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9716 (.out1(R9717), .clock(clock), .in1(R9716));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9898 (.out1(R9899), .clock(clock), .in1(R9898));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10025 (.out1(R10026), .clock(clock), .in1(R10025));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10147 (.out1(R10148), .clock(clock), .in1(R10147));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10316 (.out1(R10317), .clock(clock), .in1(R10316));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10429 (.out1(R10430), .clock(clock), .in1(R10429));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10537 (.out1(R10538), .clock(clock), .in1(R10537));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10693 (.out1(R10694), .clock(clock), .in1(R10693));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10793 (.out1(R10794), .clock(clock), .in1(R10793));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10888 (.out1(R10889), .clock(clock), .in1(R10888));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11030 (.out1(R11031), .clock(clock), .in1(R11030));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11117 (.out1(R11118), .clock(clock), .in1(R11117));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11199 (.out1(R11200), .clock(clock), .in1(R11199));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11328 (.out1(R11329), .clock(clock), .in1(R11328));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11402 (.out1(R11403), .clock(clock), .in1(off_3643));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11471 (.out1(R11472), .clock(clock), .in1(_1251));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op1294 (.out1(_1252), .in1(R11472), .in2(1 'd 1));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op1295 (.out1(ifout1295), .in1(_1252), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1363 (.out1(_1320), .in1(R11329));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1356 (.out1(_1313), .in1(R11329));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1345 (.out1(_1302), .in1(R11329));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1325 (.out1(_1282), .in1(R11329));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1364 (.out1(_1321), .in1(_1320), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1357 (.out1(_1314), .in1(_1313), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1346 (.out1(_1303), .in1(_1302), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1326 (.out1(_1283), .in1(_1282), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3864 (.out1(R3865), .clock(clock), .in1(R3864));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4120 (.out1(R4121), .clock(clock), .in1(R4120));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4375 (.out1(R4376), .clock(clock), .in1(R4375));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4620 (.out1(R4621), .clock(clock), .in1(R4620));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4860 (.out1(R4861), .clock(clock), .in1(R4860));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5147 (.out1(R5148), .clock(clock), .in1(R5147));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5379 (.out1(R5380), .clock(clock), .in1(R5379));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5606 (.out1(R5607), .clock(clock), .in1(R5606));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5880 (.out1(R5881), .clock(clock), .in1(R5880));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6098 (.out1(R6099), .clock(clock), .in1(R6098));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6311 (.out1(R6312), .clock(clock), .in1(R6311));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6572 (.out1(R6573), .clock(clock), .in1(R6572));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6777 (.out1(R6778), .clock(clock), .in1(R6777));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6977 (.out1(R6978), .clock(clock), .in1(R6977));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7224 (.out1(R7225), .clock(clock), .in1(R7224));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7416 (.out1(R7417), .clock(clock), .in1(R7416));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7603 (.out1(R7604), .clock(clock), .in1(R7603));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7837 (.out1(R7838), .clock(clock), .in1(R7837));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8016 (.out1(R8017), .clock(clock), .in1(R8016));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8190 (.out1(R8191), .clock(clock), .in1(R8190));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8411 (.out1(R8412), .clock(clock), .in1(R8411));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8577 (.out1(R8578), .clock(clock), .in1(R8577));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8738 (.out1(R8739), .clock(clock), .in1(R8738));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8946 (.out1(R8947), .clock(clock), .in1(R8946));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9099 (.out1(R9100), .clock(clock), .in1(R9099));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9247 (.out1(R9248), .clock(clock), .in1(R9247));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9442 (.out1(R9443), .clock(clock), .in1(R9442));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9582 (.out1(R9583), .clock(clock), .in1(R9582));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9717 (.out1(R9718), .clock(clock), .in1(R9717));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9899 (.out1(R9900), .clock(clock), .in1(R9899));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10026 (.out1(R10027), .clock(clock), .in1(R10026));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10148 (.out1(R10149), .clock(clock), .in1(R10148));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10317 (.out1(R10318), .clock(clock), .in1(R10317));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10430 (.out1(R10431), .clock(clock), .in1(R10430));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10538 (.out1(R10539), .clock(clock), .in1(R10538));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10694 (.out1(R10695), .clock(clock), .in1(R10694));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10794 (.out1(R10795), .clock(clock), .in1(R10794));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10889 (.out1(R10890), .clock(clock), .in1(R10889));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11031 (.out1(R11032), .clock(clock), .in1(R11031));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11118 (.out1(R11119), .clock(clock), .in1(R11118));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11200 (.out1(R11201), .clock(clock), .in1(R11200));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11329 (.out1(R11330), .clock(clock), .in1(R11329));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11403 (.out1(R11404), .clock(clock), .in1(R11403));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11472 (.out1(R11473), .clock(clock), .in1(ifout1295));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11548 (.out1(R11549), .clock(clock), .in1(_1321));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11549 (.out1(R11550), .clock(clock), .in1(_1314));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11550 (.out1(R11551), .clock(clock), .in1(_1303));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11551 (.out1(R11552), .clock(clock), .in1(_1283));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1338 (.out1(_1295), .in1(R11330));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1318 (.out1(_1275), .in1(R11330));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1307 (.out1(_1264), .in1(R11330));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1300 (.out1(_1257), .in1(R11330));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1367 (.out1(_1324), .in1(2 'd 2), .in2(R11404));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1339 (.out1(_1296), .in1(_1295), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1319 (.out1(_1276), .in1(_1275), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1308 (.out1(_1265), .in1(_1264), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1301 (.out1(_1258), .in1(_1257), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1365 (.out1(_1322), .in1(vec94_3644_D), .in2(R11549));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1358 (.out1(_1315), .in1(vec94_3644_D), .in2(R11550));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1347 (.out1(_1304), .in1(vec94_3644_D), .in2(R11551));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1327 (.out1(_1284), .in1(vec94_3644_D), .in2(R11552));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3865 (.out1(R3866), .clock(clock), .in1(R3865));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4121 (.out1(R4122), .clock(clock), .in1(R4121));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4376 (.out1(R4377), .clock(clock), .in1(R4376));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4621 (.out1(R4622), .clock(clock), .in1(R4621));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4861 (.out1(R4862), .clock(clock), .in1(R4861));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5148 (.out1(R5149), .clock(clock), .in1(R5148));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5380 (.out1(R5381), .clock(clock), .in1(R5380));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5607 (.out1(R5608), .clock(clock), .in1(R5607));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5881 (.out1(R5882), .clock(clock), .in1(R5881));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6099 (.out1(R6100), .clock(clock), .in1(R6099));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6312 (.out1(R6313), .clock(clock), .in1(R6312));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6573 (.out1(R6574), .clock(clock), .in1(R6573));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6778 (.out1(R6779), .clock(clock), .in1(R6778));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6978 (.out1(R6979), .clock(clock), .in1(R6978));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7225 (.out1(R7226), .clock(clock), .in1(R7225));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7417 (.out1(R7418), .clock(clock), .in1(R7417));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7604 (.out1(R7605), .clock(clock), .in1(R7604));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7838 (.out1(R7839), .clock(clock), .in1(R7838));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8017 (.out1(R8018), .clock(clock), .in1(R8017));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8191 (.out1(R8192), .clock(clock), .in1(R8191));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8412 (.out1(R8413), .clock(clock), .in1(R8412));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8578 (.out1(R8579), .clock(clock), .in1(R8578));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8739 (.out1(R8740), .clock(clock), .in1(R8739));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8947 (.out1(R8948), .clock(clock), .in1(R8947));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9100 (.out1(R9101), .clock(clock), .in1(R9100));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9248 (.out1(R9249), .clock(clock), .in1(R9248));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9443 (.out1(R9444), .clock(clock), .in1(R9443));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9583 (.out1(R9584), .clock(clock), .in1(R9583));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9718 (.out1(R9719), .clock(clock), .in1(R9718));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9900 (.out1(R9901), .clock(clock), .in1(R9900));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10027 (.out1(R10028), .clock(clock), .in1(R10027));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10149 (.out1(R10150), .clock(clock), .in1(R10149));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10318 (.out1(R10319), .clock(clock), .in1(R10318));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10431 (.out1(R10432), .clock(clock), .in1(R10431));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10539 (.out1(R10540), .clock(clock), .in1(R10539));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10695 (.out1(R10696), .clock(clock), .in1(R10695));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10795 (.out1(R10796), .clock(clock), .in1(R10795));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10890 (.out1(R10891), .clock(clock), .in1(R10890));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11032 (.out1(R11033), .clock(clock), .in1(R11032));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11119 (.out1(R11120), .clock(clock), .in1(R11119));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11201 (.out1(R11202), .clock(clock), .in1(R11201));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11330 (.out1(R11331), .clock(clock), .in1(R11330));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11404 (.out1(R11405), .clock(clock), .in1(R11404));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11473 (.out1(R11474), .clock(clock), .in1(R11473));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11552 (.out1(R11553), .clock(clock), .in1(_1324));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11553 (.out1(R11554), .clock(clock), .in1(_1296));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11554 (.out1(R11555), .clock(clock), .in1(_1276));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11555 (.out1(R11556), .clock(clock), .in1(_1265));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11556 (.out1(R11557), .clock(clock), .in1(_1258));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11557 (.out1(R11558), .clock(clock), .in1(_1322));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11558 (.out1(R11559), .clock(clock), .in1(_1315));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11559 (.out1(R11560), .clock(clock), .in1(_1304));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11560 (.out1(R11561), .clock(clock), .in1(_1284));
  SRAM op1366 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1323),.ADR(R11558));
  SRAM op1359 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1316),.ADR(R11559));
  SRAM op1348 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1305),.ADR(R11560));
  SRAM op1328 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1285),.ADR(R11561));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1360 (.out1(_1317), .in1(2 'd 2), .in2(R11405));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1349 (.out1(_1306), .in1(2 'd 2), .in2(R11405));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1342 (.out1(_1299), .in1(2 'd 2), .in2(R11405));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1329 (.out1(_1286), .in1(2 'd 2), .in2(R11405));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1322 (.out1(_1279), .in1(2 'd 2), .in2(R11405));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1311 (.out1(_1268), .in1(2 'd 2), .in2(R11405));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1340 (.out1(_1297), .in1(vec94_3644_D), .in2(R11554));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1320 (.out1(_1277), .in1(vec94_3644_D), .in2(R11555));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1309 (.out1(_1266), .in1(vec94_3644_D), .in2(R11556));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1302 (.out1(_1259), .in1(vec94_3644_D), .in2(R11557));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1368 (.out1(_1325), .in1(R11553), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3866 (.out1(R3867), .clock(clock), .in1(R3866));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4122 (.out1(R4123), .clock(clock), .in1(R4122));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4377 (.out1(R4378), .clock(clock), .in1(R4377));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4622 (.out1(R4623), .clock(clock), .in1(R4622));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4862 (.out1(R4863), .clock(clock), .in1(R4862));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5149 (.out1(R5150), .clock(clock), .in1(R5149));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5381 (.out1(R5382), .clock(clock), .in1(R5381));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5608 (.out1(R5609), .clock(clock), .in1(R5608));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5882 (.out1(R5883), .clock(clock), .in1(R5882));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6100 (.out1(R6101), .clock(clock), .in1(R6100));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6313 (.out1(R6314), .clock(clock), .in1(R6313));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6574 (.out1(R6575), .clock(clock), .in1(R6574));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6779 (.out1(R6780), .clock(clock), .in1(R6779));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6979 (.out1(R6980), .clock(clock), .in1(R6979));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7226 (.out1(R7227), .clock(clock), .in1(R7226));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7418 (.out1(R7419), .clock(clock), .in1(R7418));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7605 (.out1(R7606), .clock(clock), .in1(R7605));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7839 (.out1(R7840), .clock(clock), .in1(R7839));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8018 (.out1(R8019), .clock(clock), .in1(R8018));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8192 (.out1(R8193), .clock(clock), .in1(R8192));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8413 (.out1(R8414), .clock(clock), .in1(R8413));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8579 (.out1(R8580), .clock(clock), .in1(R8579));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8740 (.out1(R8741), .clock(clock), .in1(R8740));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8948 (.out1(R8949), .clock(clock), .in1(R8948));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9101 (.out1(R9102), .clock(clock), .in1(R9101));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9249 (.out1(R9250), .clock(clock), .in1(R9249));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9444 (.out1(R9445), .clock(clock), .in1(R9444));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9584 (.out1(R9585), .clock(clock), .in1(R9584));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9719 (.out1(R9720), .clock(clock), .in1(R9719));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9901 (.out1(R9902), .clock(clock), .in1(R9901));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10028 (.out1(R10029), .clock(clock), .in1(R10028));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10150 (.out1(R10151), .clock(clock), .in1(R10150));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10319 (.out1(R10320), .clock(clock), .in1(R10319));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10432 (.out1(R10433), .clock(clock), .in1(R10432));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10540 (.out1(R10541), .clock(clock), .in1(R10540));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10696 (.out1(R10697), .clock(clock), .in1(R10696));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10796 (.out1(R10797), .clock(clock), .in1(R10796));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10891 (.out1(R10892), .clock(clock), .in1(R10891));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11033 (.out1(R11034), .clock(clock), .in1(R11033));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11120 (.out1(R11121), .clock(clock), .in1(R11120));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11202 (.out1(R11203), .clock(clock), .in1(R11202));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11331 (.out1(R11332), .clock(clock), .in1(R11331));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11405 (.out1(R11406), .clock(clock), .in1(R11405));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11474 (.out1(R11475), .clock(clock), .in1(R11474));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11561 (.out1(R11562), .clock(clock), .in1(_1323));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11562 (.out1(R11563), .clock(clock), .in1(_1316));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11563 (.out1(R11564), .clock(clock), .in1(_1305));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11564 (.out1(R11565), .clock(clock), .in1(_1285));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11565 (.out1(R11566), .clock(clock), .in1(_1317));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11566 (.out1(R11567), .clock(clock), .in1(_1306));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11567 (.out1(R11568), .clock(clock), .in1(_1299));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11568 (.out1(R11569), .clock(clock), .in1(_1286));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11569 (.out1(R11570), .clock(clock), .in1(_1279));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11570 (.out1(R11571), .clock(clock), .in1(_1268));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11571 (.out1(R11572), .clock(clock), .in1(_1297));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11572 (.out1(R11573), .clock(clock), .in1(_1277));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11573 (.out1(R11574), .clock(clock), .in1(_1266));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11574 (.out1(R11575), .clock(clock), .in1(_1259));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11575 (.out1(R11576), .clock(clock), .in1(_1325));
  SRAM op1341 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1298),.ADR(R11572));
  SRAM op1321 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1278),.ADR(R11573));
  SRAM op1310 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1267),.ADR(R11574));
  SRAM op1303 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1260),.ADR(R11575));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1369 (.out1(_1326), .in1(R11562), .in2(R11576));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1370 (.out1(_1327), .in1(_1326), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1361 (.out1(_1318), .in1(R11566), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1350 (.out1(_1307), .in1(R11567), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1330 (.out1(_1287), .in1(R11569), .in2(64 'd 18446744073709551615));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1304 (.out1(_1261), .in1(2 'd 2), .in2(R11406));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1371 (.out1(_1328), .in1(_1327), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1362 (.out1(_1319), .in1(R11563), .in2(_1318));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1351 (.out1(_1308), .in1(R11564), .in2(_1307));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1331 (.out1(_1288), .in1(R11565), .in2(_1287));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1372 (.out1(_1329), .in1(_1319), .in2(_1328));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1352 (.out1(_1309), .in1(_1308), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1343 (.out1(_1300), .in1(R11568), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1332 (.out1(_1289), .in1(_1288), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1323 (.out1(_1280), .in1(R11570), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1312 (.out1(_1269), .in1(R11571), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3867 (.out1(R3868), .clock(clock), .in1(R3867));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4123 (.out1(R4124), .clock(clock), .in1(R4123));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4378 (.out1(R4379), .clock(clock), .in1(R4378));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4623 (.out1(R4624), .clock(clock), .in1(R4623));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4863 (.out1(R4864), .clock(clock), .in1(R4863));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5150 (.out1(R5151), .clock(clock), .in1(R5150));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5382 (.out1(R5383), .clock(clock), .in1(R5382));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5609 (.out1(R5610), .clock(clock), .in1(R5609));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5883 (.out1(R5884), .clock(clock), .in1(R5883));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6101 (.out1(R6102), .clock(clock), .in1(R6101));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6314 (.out1(R6315), .clock(clock), .in1(R6314));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6575 (.out1(R6576), .clock(clock), .in1(R6575));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6780 (.out1(R6781), .clock(clock), .in1(R6780));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6980 (.out1(R6981), .clock(clock), .in1(R6980));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7227 (.out1(R7228), .clock(clock), .in1(R7227));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7419 (.out1(R7420), .clock(clock), .in1(R7419));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7606 (.out1(R7607), .clock(clock), .in1(R7606));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7840 (.out1(R7841), .clock(clock), .in1(R7840));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8019 (.out1(R8020), .clock(clock), .in1(R8019));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8193 (.out1(R8194), .clock(clock), .in1(R8193));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8414 (.out1(R8415), .clock(clock), .in1(R8414));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8580 (.out1(R8581), .clock(clock), .in1(R8580));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8741 (.out1(R8742), .clock(clock), .in1(R8741));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8949 (.out1(R8950), .clock(clock), .in1(R8949));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9102 (.out1(R9103), .clock(clock), .in1(R9102));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9250 (.out1(R9251), .clock(clock), .in1(R9250));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9445 (.out1(R9446), .clock(clock), .in1(R9445));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9585 (.out1(R9586), .clock(clock), .in1(R9585));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9720 (.out1(R9721), .clock(clock), .in1(R9720));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9902 (.out1(R9903), .clock(clock), .in1(R9902));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10029 (.out1(R10030), .clock(clock), .in1(R10029));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10151 (.out1(R10152), .clock(clock), .in1(R10151));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10320 (.out1(R10321), .clock(clock), .in1(R10320));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10433 (.out1(R10434), .clock(clock), .in1(R10433));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10541 (.out1(R10542), .clock(clock), .in1(R10541));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10697 (.out1(R10698), .clock(clock), .in1(R10697));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10797 (.out1(R10798), .clock(clock), .in1(R10797));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10892 (.out1(R10893), .clock(clock), .in1(R10892));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11034 (.out1(R11035), .clock(clock), .in1(R11034));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11121 (.out1(R11122), .clock(clock), .in1(R11121));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11203 (.out1(R11204), .clock(clock), .in1(R11203));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11332 (.out1(R11333), .clock(clock), .in1(R11332));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11406 (.out1(R11407), .clock(clock), .in1(R11406));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11475 (.out1(R11476), .clock(clock), .in1(R11475));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11576 (.out1(R11577), .clock(clock), .in1(_1298));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11577 (.out1(R11578), .clock(clock), .in1(_1278));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11578 (.out1(R11579), .clock(clock), .in1(_1267));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11579 (.out1(R11580), .clock(clock), .in1(_1260));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11580 (.out1(R11581), .clock(clock), .in1(_1261));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11581 (.out1(R11582), .clock(clock), .in1(_1329));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11582 (.out1(R11583), .clock(clock), .in1(_1309));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11583 (.out1(R11584), .clock(clock), .in1(_1300));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11584 (.out1(R11585), .clock(clock), .in1(_1289));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11585 (.out1(R11586), .clock(clock), .in1(_1280));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11586 (.out1(R11587), .clock(clock), .in1(_1269));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1353 (.out1(_1310), .in1(R11583), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1344 (.out1(_1301), .in1(R11577), .in2(R11584));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1313 (.out1(_1270), .in1(R11579), .in2(R11587));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1373 (.out1(_1330), .in1(R11582), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1354 (.out1(_1311), .in1(_1301), .in2(_1310));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1333 (.out1(_1290), .in1(R11585), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1324 (.out1(_1281), .in1(R11578), .in2(R11586));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1314 (.out1(_1271), .in1(_1270), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1305 (.out1(_1262), .in1(R11581), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1334 (.out1(_1291), .in1(_1281), .in2(_1290));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1374 (.out1(_1331), .in1(_1330), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1355 (.out1(_1312), .in1(_1311), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1315 (.out1(_1272), .in1(_1271), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1306 (.out1(_1263), .in1(R11580), .in2(_1262));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1375 (.out1(_1332), .in1(_1312), .in2(_1331));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1335 (.out1(_1292), .in1(_1291), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1316 (.out1(_1273), .in1(_1263), .in2(_1272));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3868 (.out1(R3869), .clock(clock), .in1(R3868));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4124 (.out1(R4125), .clock(clock), .in1(R4124));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4379 (.out1(R4380), .clock(clock), .in1(R4379));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4624 (.out1(R4625), .clock(clock), .in1(R4624));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4864 (.out1(R4865), .clock(clock), .in1(R4864));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5151 (.out1(R5152), .clock(clock), .in1(R5151));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5383 (.out1(R5384), .clock(clock), .in1(R5383));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5610 (.out1(R5611), .clock(clock), .in1(R5610));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5884 (.out1(R5885), .clock(clock), .in1(R5884));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6102 (.out1(R6103), .clock(clock), .in1(R6102));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6315 (.out1(R6316), .clock(clock), .in1(R6315));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6576 (.out1(R6577), .clock(clock), .in1(R6576));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6781 (.out1(R6782), .clock(clock), .in1(R6781));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6981 (.out1(R6982), .clock(clock), .in1(R6981));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7228 (.out1(R7229), .clock(clock), .in1(R7228));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7420 (.out1(R7421), .clock(clock), .in1(R7420));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7607 (.out1(R7608), .clock(clock), .in1(R7607));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7841 (.out1(R7842), .clock(clock), .in1(R7841));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8020 (.out1(R8021), .clock(clock), .in1(R8020));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8194 (.out1(R8195), .clock(clock), .in1(R8194));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8415 (.out1(R8416), .clock(clock), .in1(R8415));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8581 (.out1(R8582), .clock(clock), .in1(R8581));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8742 (.out1(R8743), .clock(clock), .in1(R8742));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8950 (.out1(R8951), .clock(clock), .in1(R8950));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9103 (.out1(R9104), .clock(clock), .in1(R9103));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9251 (.out1(R9252), .clock(clock), .in1(R9251));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9446 (.out1(R9447), .clock(clock), .in1(R9446));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9586 (.out1(R9587), .clock(clock), .in1(R9586));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9721 (.out1(R9722), .clock(clock), .in1(R9721));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9903 (.out1(R9904), .clock(clock), .in1(R9903));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10030 (.out1(R10031), .clock(clock), .in1(R10030));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10152 (.out1(R10153), .clock(clock), .in1(R10152));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10321 (.out1(R10322), .clock(clock), .in1(R10321));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10434 (.out1(R10435), .clock(clock), .in1(R10434));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10542 (.out1(R10543), .clock(clock), .in1(R10542));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10698 (.out1(R10699), .clock(clock), .in1(R10698));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10798 (.out1(R10799), .clock(clock), .in1(R10798));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10893 (.out1(R10894), .clock(clock), .in1(R10893));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11035 (.out1(R11036), .clock(clock), .in1(R11035));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11122 (.out1(R11123), .clock(clock), .in1(R11122));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11204 (.out1(R11205), .clock(clock), .in1(R11204));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11333 (.out1(R11334), .clock(clock), .in1(R11333));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11407 (.out1(R11408), .clock(clock), .in1(R11407));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11476 (.out1(R11477), .clock(clock), .in1(R11476));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11587 (.out1(R11588), .clock(clock), .in1(_1332));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11588 (.out1(R11589), .clock(clock), .in1(_1292));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11589 (.out1(R11590), .clock(clock), .in1(_1273));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1296 (.out1(_1253), .in1(R11334));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1336 (.out1(_1293), .in1(R11589), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1317 (.out1(_1274), .in1(R11590), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op1376 (.out1(_1333), .in1(R11588), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1337 (.out1(_1294), .in1(_1274), .in2(_1293));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1297 (.out1(_1254), .in1(_1253), .in2(2 'd 2));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1377 (.out1(_1334), .in1(_1294), .in2(_1333));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op1378 (.out1(_1335), .in1(_1334), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3869 (.out1(R3870), .clock(clock), .in1(R3869));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4125 (.out1(R4126), .clock(clock), .in1(R4125));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4380 (.out1(R4381), .clock(clock), .in1(R4380));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4625 (.out1(R4626), .clock(clock), .in1(R4625));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4865 (.out1(R4866), .clock(clock), .in1(R4865));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5152 (.out1(R5153), .clock(clock), .in1(R5152));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5384 (.out1(R5385), .clock(clock), .in1(R5384));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5611 (.out1(R5612), .clock(clock), .in1(R5611));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5885 (.out1(R5886), .clock(clock), .in1(R5885));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6103 (.out1(R6104), .clock(clock), .in1(R6103));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6316 (.out1(R6317), .clock(clock), .in1(R6316));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6577 (.out1(R6578), .clock(clock), .in1(R6577));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6782 (.out1(R6783), .clock(clock), .in1(R6782));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6982 (.out1(R6983), .clock(clock), .in1(R6982));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7229 (.out1(R7230), .clock(clock), .in1(R7229));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7421 (.out1(R7422), .clock(clock), .in1(R7421));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7608 (.out1(R7609), .clock(clock), .in1(R7608));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7842 (.out1(R7843), .clock(clock), .in1(R7842));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8021 (.out1(R8022), .clock(clock), .in1(R8021));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8195 (.out1(R8196), .clock(clock), .in1(R8195));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8416 (.out1(R8417), .clock(clock), .in1(R8416));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8582 (.out1(R8583), .clock(clock), .in1(R8582));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8743 (.out1(R8744), .clock(clock), .in1(R8743));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8951 (.out1(R8952), .clock(clock), .in1(R8951));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9104 (.out1(R9105), .clock(clock), .in1(R9104));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9252 (.out1(R9253), .clock(clock), .in1(R9252));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9447 (.out1(R9448), .clock(clock), .in1(R9447));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9587 (.out1(R9588), .clock(clock), .in1(R9587));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9722 (.out1(R9723), .clock(clock), .in1(R9722));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9904 (.out1(R9905), .clock(clock), .in1(R9904));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10031 (.out1(R10032), .clock(clock), .in1(R10031));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10153 (.out1(R10154), .clock(clock), .in1(R10153));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10322 (.out1(R10323), .clock(clock), .in1(R10322));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10435 (.out1(R10436), .clock(clock), .in1(R10435));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10543 (.out1(R10544), .clock(clock), .in1(R10543));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10699 (.out1(R10700), .clock(clock), .in1(R10699));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10799 (.out1(R10800), .clock(clock), .in1(R10799));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10894 (.out1(R10895), .clock(clock), .in1(R10894));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11036 (.out1(R11037), .clock(clock), .in1(R11036));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11123 (.out1(R11124), .clock(clock), .in1(R11123));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11205 (.out1(R11206), .clock(clock), .in1(R11205));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11334 (.out1(R11335), .clock(clock), .in1(R11334));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11408 (.out1(R11409), .clock(clock), .in1(R11408));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11477 (.out1(R11478), .clock(clock), .in1(R11477));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11590 (.out1(R11591), .clock(clock), .in1(_1254));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11591 (.out1(R11592), .clock(clock), .in1(_1335));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op1379 (.out1(_1336), .in1(R11592), .in2(57 'd 72340172838076673));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1298 (.out1(_1255), .in1(base0_94_3649_D), .in2(R11591));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3870 (.out1(R3871), .clock(clock), .in1(R3870));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4126 (.out1(R4127), .clock(clock), .in1(R4126));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4381 (.out1(R4382), .clock(clock), .in1(R4381));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4626 (.out1(R4627), .clock(clock), .in1(R4626));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4866 (.out1(R4867), .clock(clock), .in1(R4866));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5153 (.out1(R5154), .clock(clock), .in1(R5153));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5385 (.out1(R5386), .clock(clock), .in1(R5385));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5612 (.out1(R5613), .clock(clock), .in1(R5612));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5886 (.out1(R5887), .clock(clock), .in1(R5886));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6104 (.out1(R6105), .clock(clock), .in1(R6104));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6317 (.out1(R6318), .clock(clock), .in1(R6317));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6578 (.out1(R6579), .clock(clock), .in1(R6578));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6783 (.out1(R6784), .clock(clock), .in1(R6783));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6983 (.out1(R6984), .clock(clock), .in1(R6983));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7230 (.out1(R7231), .clock(clock), .in1(R7230));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7422 (.out1(R7423), .clock(clock), .in1(R7422));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7609 (.out1(R7610), .clock(clock), .in1(R7609));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7843 (.out1(R7844), .clock(clock), .in1(R7843));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8022 (.out1(R8023), .clock(clock), .in1(R8022));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8196 (.out1(R8197), .clock(clock), .in1(R8196));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8417 (.out1(R8418), .clock(clock), .in1(R8417));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8583 (.out1(R8584), .clock(clock), .in1(R8583));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8744 (.out1(R8745), .clock(clock), .in1(R8744));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8952 (.out1(R8953), .clock(clock), .in1(R8952));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9105 (.out1(R9106), .clock(clock), .in1(R9105));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9253 (.out1(R9254), .clock(clock), .in1(R9253));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9448 (.out1(R9449), .clock(clock), .in1(R9448));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9588 (.out1(R9589), .clock(clock), .in1(R9588));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9723 (.out1(R9724), .clock(clock), .in1(R9723));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9905 (.out1(R9906), .clock(clock), .in1(R9905));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10032 (.out1(R10033), .clock(clock), .in1(R10032));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10154 (.out1(R10155), .clock(clock), .in1(R10154));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10323 (.out1(R10324), .clock(clock), .in1(R10323));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10436 (.out1(R10437), .clock(clock), .in1(R10436));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10544 (.out1(R10545), .clock(clock), .in1(R10544));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10700 (.out1(R10701), .clock(clock), .in1(R10700));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10800 (.out1(R10801), .clock(clock), .in1(R10800));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10895 (.out1(R10896), .clock(clock), .in1(R10895));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11037 (.out1(R11038), .clock(clock), .in1(R11037));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11124 (.out1(R11125), .clock(clock), .in1(R11124));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11206 (.out1(R11207), .clock(clock), .in1(R11206));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11335 (.out1(R11336), .clock(clock), .in1(R11335));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11409 (.out1(R11410), .clock(clock), .in1(R11409));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11478 (.out1(R11479), .clock(clock), .in1(R11478));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11592 (.out1(R11593), .clock(clock), .in1(_1336));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11593 (.out1(R11594), .clock(clock), .in1(_1255));
  SRAM op1299 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1256),.ADR(R11594));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op1380 (.out1(_1337), .in1(R11593), .in2(6 'd 56));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3871 (.out1(R3872), .clock(clock), .in1(R3871));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4127 (.out1(R4128), .clock(clock), .in1(R4127));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4382 (.out1(R4383), .clock(clock), .in1(R4382));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4627 (.out1(R4628), .clock(clock), .in1(R4627));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4867 (.out1(R4868), .clock(clock), .in1(R4867));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5154 (.out1(R5155), .clock(clock), .in1(R5154));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5386 (.out1(R5387), .clock(clock), .in1(R5386));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5613 (.out1(R5614), .clock(clock), .in1(R5613));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5887 (.out1(R5888), .clock(clock), .in1(R5887));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6105 (.out1(R6106), .clock(clock), .in1(R6105));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6318 (.out1(R6319), .clock(clock), .in1(R6318));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6579 (.out1(R6580), .clock(clock), .in1(R6579));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6784 (.out1(R6785), .clock(clock), .in1(R6784));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6984 (.out1(R6985), .clock(clock), .in1(R6984));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7231 (.out1(R7232), .clock(clock), .in1(R7231));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7423 (.out1(R7424), .clock(clock), .in1(R7423));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7610 (.out1(R7611), .clock(clock), .in1(R7610));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7844 (.out1(R7845), .clock(clock), .in1(R7844));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8023 (.out1(R8024), .clock(clock), .in1(R8023));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8197 (.out1(R8198), .clock(clock), .in1(R8197));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8418 (.out1(R8419), .clock(clock), .in1(R8418));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8584 (.out1(R8585), .clock(clock), .in1(R8584));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8745 (.out1(R8746), .clock(clock), .in1(R8745));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8953 (.out1(R8954), .clock(clock), .in1(R8953));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9106 (.out1(R9107), .clock(clock), .in1(R9106));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9254 (.out1(R9255), .clock(clock), .in1(R9254));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9449 (.out1(R9450), .clock(clock), .in1(R9449));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9589 (.out1(R9590), .clock(clock), .in1(R9589));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9724 (.out1(R9725), .clock(clock), .in1(R9724));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9906 (.out1(R9907), .clock(clock), .in1(R9906));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10033 (.out1(R10034), .clock(clock), .in1(R10033));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10155 (.out1(R10156), .clock(clock), .in1(R10155));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10324 (.out1(R10325), .clock(clock), .in1(R10324));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10437 (.out1(R10438), .clock(clock), .in1(R10437));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10545 (.out1(R10546), .clock(clock), .in1(R10545));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10701 (.out1(R10702), .clock(clock), .in1(R10701));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10801 (.out1(R10802), .clock(clock), .in1(R10801));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10896 (.out1(R10897), .clock(clock), .in1(R10896));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11038 (.out1(R11039), .clock(clock), .in1(R11038));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11125 (.out1(R11126), .clock(clock), .in1(R11125));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11207 (.out1(R11208), .clock(clock), .in1(R11207));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11336 (.out1(R11337), .clock(clock), .in1(R11336));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11410 (.out1(R11411), .clock(clock), .in1(R11410));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11479 (.out1(R11480), .clock(clock), .in1(R11479));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11594 (.out1(R11595), .clock(clock), .in1(_1256));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11595 (.out1(R11596), .clock(clock), .in1(_1337));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1381 (.out1(_1338), .in1(R11596));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1382 (.out1(_1339), .in1(R11595), .in2(_1338));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1383 (.out1(idx_3650), .in1(_1339), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3872 (.out1(R3873), .clock(clock), .in1(R3872));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4128 (.out1(R4129), .clock(clock), .in1(R4128));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4383 (.out1(R4384), .clock(clock), .in1(R4383));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4628 (.out1(R4629), .clock(clock), .in1(R4628));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4868 (.out1(R4869), .clock(clock), .in1(R4868));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5155 (.out1(R5156), .clock(clock), .in1(R5155));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5387 (.out1(R5388), .clock(clock), .in1(R5387));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5614 (.out1(R5615), .clock(clock), .in1(R5614));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5888 (.out1(R5889), .clock(clock), .in1(R5888));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6106 (.out1(R6107), .clock(clock), .in1(R6106));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6319 (.out1(R6320), .clock(clock), .in1(R6319));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6580 (.out1(R6581), .clock(clock), .in1(R6580));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6785 (.out1(R6786), .clock(clock), .in1(R6785));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6985 (.out1(R6986), .clock(clock), .in1(R6985));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7232 (.out1(R7233), .clock(clock), .in1(R7232));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7424 (.out1(R7425), .clock(clock), .in1(R7424));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7611 (.out1(R7612), .clock(clock), .in1(R7611));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7845 (.out1(R7846), .clock(clock), .in1(R7845));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8024 (.out1(R8025), .clock(clock), .in1(R8024));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8198 (.out1(R8199), .clock(clock), .in1(R8198));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8419 (.out1(R8420), .clock(clock), .in1(R8419));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8585 (.out1(R8586), .clock(clock), .in1(R8585));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8746 (.out1(R8747), .clock(clock), .in1(R8746));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8954 (.out1(R8955), .clock(clock), .in1(R8954));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9107 (.out1(R9108), .clock(clock), .in1(R9107));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9255 (.out1(R9256), .clock(clock), .in1(R9255));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9450 (.out1(R9451), .clock(clock), .in1(R9450));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9590 (.out1(R9591), .clock(clock), .in1(R9590));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9725 (.out1(R9726), .clock(clock), .in1(R9725));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9907 (.out1(R9908), .clock(clock), .in1(R9907));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10034 (.out1(R10035), .clock(clock), .in1(R10034));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10156 (.out1(R10157), .clock(clock), .in1(R10156));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10325 (.out1(R10326), .clock(clock), .in1(R10325));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10438 (.out1(R10439), .clock(clock), .in1(R10438));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10546 (.out1(R10547), .clock(clock), .in1(R10546));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10702 (.out1(R10703), .clock(clock), .in1(R10702));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10802 (.out1(R10803), .clock(clock), .in1(R10802));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10897 (.out1(R10898), .clock(clock), .in1(R10897));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11039 (.out1(R11040), .clock(clock), .in1(R11039));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11126 (.out1(R11127), .clock(clock), .in1(R11126));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11208 (.out1(R11209), .clock(clock), .in1(R11208));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11337 (.out1(R11338), .clock(clock), .in1(R11337));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11411 (.out1(R11412), .clock(clock), .in1(R11411));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11480 (.out1(R11481), .clock(clock), .in1(R11480));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11596 (.out1(R11597), .clock(clock), .in1(idx_3650));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1387 (.out1(_1342), .in1(R11597));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1388 (.out1(_1343), .in1(_1342), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3873 (.out1(R3874), .clock(clock), .in1(R3873));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4129 (.out1(R4130), .clock(clock), .in1(R4129));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4384 (.out1(R4385), .clock(clock), .in1(R4384));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4629 (.out1(R4630), .clock(clock), .in1(R4629));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4869 (.out1(R4870), .clock(clock), .in1(R4869));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5156 (.out1(R5157), .clock(clock), .in1(R5156));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5388 (.out1(R5389), .clock(clock), .in1(R5388));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5615 (.out1(R5616), .clock(clock), .in1(R5615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5889 (.out1(R5890), .clock(clock), .in1(R5889));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6107 (.out1(R6108), .clock(clock), .in1(R6107));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6320 (.out1(R6321), .clock(clock), .in1(R6320));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6581 (.out1(R6582), .clock(clock), .in1(R6581));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6786 (.out1(R6787), .clock(clock), .in1(R6786));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6986 (.out1(R6987), .clock(clock), .in1(R6986));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7233 (.out1(R7234), .clock(clock), .in1(R7233));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7425 (.out1(R7426), .clock(clock), .in1(R7425));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7612 (.out1(R7613), .clock(clock), .in1(R7612));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7846 (.out1(R7847), .clock(clock), .in1(R7846));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8025 (.out1(R8026), .clock(clock), .in1(R8025));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8199 (.out1(R8200), .clock(clock), .in1(R8199));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8420 (.out1(R8421), .clock(clock), .in1(R8420));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8586 (.out1(R8587), .clock(clock), .in1(R8586));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8747 (.out1(R8748), .clock(clock), .in1(R8747));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8955 (.out1(R8956), .clock(clock), .in1(R8955));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9108 (.out1(R9109), .clock(clock), .in1(R9108));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9256 (.out1(R9257), .clock(clock), .in1(R9256));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9451 (.out1(R9452), .clock(clock), .in1(R9451));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9591 (.out1(R9592), .clock(clock), .in1(R9591));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9726 (.out1(R9727), .clock(clock), .in1(R9726));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9908 (.out1(R9909), .clock(clock), .in1(R9908));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10035 (.out1(R10036), .clock(clock), .in1(R10035));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10157 (.out1(R10158), .clock(clock), .in1(R10157));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10326 (.out1(R10327), .clock(clock), .in1(R10326));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10439 (.out1(R10440), .clock(clock), .in1(R10439));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10547 (.out1(R10548), .clock(clock), .in1(R10547));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10703 (.out1(R10704), .clock(clock), .in1(R10703));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10803 (.out1(R10804), .clock(clock), .in1(R10803));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10898 (.out1(R10899), .clock(clock), .in1(R10898));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11040 (.out1(R11041), .clock(clock), .in1(R11040));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11127 (.out1(R11128), .clock(clock), .in1(R11127));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11209 (.out1(R11210), .clock(clock), .in1(R11209));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11338 (.out1(R11339), .clock(clock), .in1(R11338));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11412 (.out1(R11413), .clock(clock), .in1(R11412));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11481 (.out1(R11482), .clock(clock), .in1(R11481));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11597 (.out1(R11598), .clock(clock), .in1(R11597));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11658 (.out1(R11659), .clock(clock), .in1(_1343));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1389 (.out1(_1344), .in1(vec100_3652_D), .in2(R11659));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3874 (.out1(R3875), .clock(clock), .in1(R3874));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4130 (.out1(R4131), .clock(clock), .in1(R4130));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4385 (.out1(R4386), .clock(clock), .in1(R4385));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4630 (.out1(R4631), .clock(clock), .in1(R4630));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4870 (.out1(R4871), .clock(clock), .in1(R4870));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5157 (.out1(R5158), .clock(clock), .in1(R5157));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5389 (.out1(R5390), .clock(clock), .in1(R5389));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5616 (.out1(R5617), .clock(clock), .in1(R5616));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5890 (.out1(R5891), .clock(clock), .in1(R5890));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6108 (.out1(R6109), .clock(clock), .in1(R6108));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6321 (.out1(R6322), .clock(clock), .in1(R6321));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6582 (.out1(R6583), .clock(clock), .in1(R6582));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6787 (.out1(R6788), .clock(clock), .in1(R6787));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6987 (.out1(R6988), .clock(clock), .in1(R6987));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7234 (.out1(R7235), .clock(clock), .in1(R7234));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7426 (.out1(R7427), .clock(clock), .in1(R7426));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7613 (.out1(R7614), .clock(clock), .in1(R7613));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7847 (.out1(R7848), .clock(clock), .in1(R7847));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8026 (.out1(R8027), .clock(clock), .in1(R8026));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8200 (.out1(R8201), .clock(clock), .in1(R8200));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8421 (.out1(R8422), .clock(clock), .in1(R8421));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8587 (.out1(R8588), .clock(clock), .in1(R8587));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8748 (.out1(R8749), .clock(clock), .in1(R8748));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8956 (.out1(R8957), .clock(clock), .in1(R8956));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9109 (.out1(R9110), .clock(clock), .in1(R9109));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9257 (.out1(R9258), .clock(clock), .in1(R9257));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9452 (.out1(R9453), .clock(clock), .in1(R9452));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9592 (.out1(R9593), .clock(clock), .in1(R9592));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9727 (.out1(R9728), .clock(clock), .in1(R9727));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9909 (.out1(R9910), .clock(clock), .in1(R9909));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10036 (.out1(R10037), .clock(clock), .in1(R10036));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10158 (.out1(R10159), .clock(clock), .in1(R10158));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10327 (.out1(R10328), .clock(clock), .in1(R10327));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10440 (.out1(R10441), .clock(clock), .in1(R10440));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10548 (.out1(R10549), .clock(clock), .in1(R10548));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10704 (.out1(R10705), .clock(clock), .in1(R10704));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10804 (.out1(R10805), .clock(clock), .in1(R10804));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10899 (.out1(R10900), .clock(clock), .in1(R10899));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11041 (.out1(R11042), .clock(clock), .in1(R11041));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11128 (.out1(R11129), .clock(clock), .in1(R11128));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11210 (.out1(R11211), .clock(clock), .in1(R11210));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11339 (.out1(R11340), .clock(clock), .in1(R11339));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11413 (.out1(R11414), .clock(clock), .in1(R11413));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11482 (.out1(R11483), .clock(clock), .in1(R11482));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11598 (.out1(R11599), .clock(clock), .in1(R11598));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11659 (.out1(R11660), .clock(clock), .in1(_1344));
  SRAM op1390 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1345),.ADR(R11660));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3875 (.out1(R3876), .clock(clock), .in1(R3875));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4131 (.out1(R4132), .clock(clock), .in1(R4131));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4386 (.out1(R4387), .clock(clock), .in1(R4386));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4631 (.out1(R4632), .clock(clock), .in1(R4631));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4871 (.out1(R4872), .clock(clock), .in1(R4871));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5158 (.out1(R5159), .clock(clock), .in1(R5158));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5390 (.out1(R5391), .clock(clock), .in1(R5390));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5617 (.out1(R5618), .clock(clock), .in1(R5617));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5891 (.out1(R5892), .clock(clock), .in1(R5891));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6109 (.out1(R6110), .clock(clock), .in1(R6109));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6322 (.out1(R6323), .clock(clock), .in1(R6322));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6583 (.out1(R6584), .clock(clock), .in1(R6583));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6788 (.out1(R6789), .clock(clock), .in1(R6788));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6988 (.out1(R6989), .clock(clock), .in1(R6988));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7235 (.out1(R7236), .clock(clock), .in1(R7235));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7427 (.out1(R7428), .clock(clock), .in1(R7427));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7614 (.out1(R7615), .clock(clock), .in1(R7614));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7848 (.out1(R7849), .clock(clock), .in1(R7848));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8027 (.out1(R8028), .clock(clock), .in1(R8027));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8201 (.out1(R8202), .clock(clock), .in1(R8201));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8422 (.out1(R8423), .clock(clock), .in1(R8422));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8588 (.out1(R8589), .clock(clock), .in1(R8588));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8749 (.out1(R8750), .clock(clock), .in1(R8749));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8957 (.out1(R8958), .clock(clock), .in1(R8957));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9110 (.out1(R9111), .clock(clock), .in1(R9110));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9258 (.out1(R9259), .clock(clock), .in1(R9258));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9453 (.out1(R9454), .clock(clock), .in1(R9453));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9593 (.out1(R9594), .clock(clock), .in1(R9593));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9728 (.out1(R9729), .clock(clock), .in1(R9728));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9910 (.out1(R9911), .clock(clock), .in1(R9910));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10037 (.out1(R10038), .clock(clock), .in1(R10037));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10159 (.out1(R10160), .clock(clock), .in1(R10159));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10328 (.out1(R10329), .clock(clock), .in1(R10328));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10441 (.out1(R10442), .clock(clock), .in1(R10441));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10549 (.out1(R10550), .clock(clock), .in1(R10549));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10705 (.out1(R10706), .clock(clock), .in1(R10705));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10805 (.out1(R10806), .clock(clock), .in1(R10805));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10900 (.out1(R10901), .clock(clock), .in1(R10900));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11042 (.out1(R11043), .clock(clock), .in1(R11042));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11129 (.out1(R11130), .clock(clock), .in1(R11129));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11211 (.out1(R11212), .clock(clock), .in1(R11211));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11340 (.out1(R11341), .clock(clock), .in1(R11340));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11414 (.out1(R11415), .clock(clock), .in1(R11414));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11483 (.out1(R11484), .clock(clock), .in1(R11483));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11599 (.out1(R11600), .clock(clock), .in1(R11599));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11660 (.out1(R11661), .clock(clock), .in1(_1345));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(5), .BITSIZE_out1(64), .PRECISION(64)) op1384 (.out1(_1340), .in1(ip2_3602_D), .in2(5 'd 22));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1385 (.out1(_1341), .in1(_1340));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op1386 (.out1(off_3651), .in1(_1341), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1391 (.out1(_1346), .in1(R11661), .in2(off_3651));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3876 (.out1(R3877), .clock(clock), .in1(R3876));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4132 (.out1(R4133), .clock(clock), .in1(R4132));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4387 (.out1(R4388), .clock(clock), .in1(R4387));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4632 (.out1(R4633), .clock(clock), .in1(R4632));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4872 (.out1(R4873), .clock(clock), .in1(R4872));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5159 (.out1(R5160), .clock(clock), .in1(R5159));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5391 (.out1(R5392), .clock(clock), .in1(R5391));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5618 (.out1(R5619), .clock(clock), .in1(R5618));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5892 (.out1(R5893), .clock(clock), .in1(R5892));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6110 (.out1(R6111), .clock(clock), .in1(R6110));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6323 (.out1(R6324), .clock(clock), .in1(R6323));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6584 (.out1(R6585), .clock(clock), .in1(R6584));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6789 (.out1(R6790), .clock(clock), .in1(R6789));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6989 (.out1(R6990), .clock(clock), .in1(R6989));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7236 (.out1(R7237), .clock(clock), .in1(R7236));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7428 (.out1(R7429), .clock(clock), .in1(R7428));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7615 (.out1(R7616), .clock(clock), .in1(R7615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7849 (.out1(R7850), .clock(clock), .in1(R7849));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8028 (.out1(R8029), .clock(clock), .in1(R8028));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8202 (.out1(R8203), .clock(clock), .in1(R8202));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8423 (.out1(R8424), .clock(clock), .in1(R8423));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8589 (.out1(R8590), .clock(clock), .in1(R8589));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8750 (.out1(R8751), .clock(clock), .in1(R8750));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8958 (.out1(R8959), .clock(clock), .in1(R8958));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9111 (.out1(R9112), .clock(clock), .in1(R9111));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9259 (.out1(R9260), .clock(clock), .in1(R9259));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9454 (.out1(R9455), .clock(clock), .in1(R9454));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9594 (.out1(R9595), .clock(clock), .in1(R9594));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9729 (.out1(R9730), .clock(clock), .in1(R9729));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9911 (.out1(R9912), .clock(clock), .in1(R9911));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10038 (.out1(R10039), .clock(clock), .in1(R10038));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10160 (.out1(R10161), .clock(clock), .in1(R10160));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10329 (.out1(R10330), .clock(clock), .in1(R10329));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10442 (.out1(R10443), .clock(clock), .in1(R10442));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10550 (.out1(R10551), .clock(clock), .in1(R10550));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10706 (.out1(R10707), .clock(clock), .in1(R10706));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10806 (.out1(R10807), .clock(clock), .in1(R10806));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10901 (.out1(R10902), .clock(clock), .in1(R10901));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11043 (.out1(R11044), .clock(clock), .in1(R11043));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11130 (.out1(R11131), .clock(clock), .in1(R11130));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11212 (.out1(R11213), .clock(clock), .in1(R11212));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11341 (.out1(R11342), .clock(clock), .in1(R11341));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11415 (.out1(R11416), .clock(clock), .in1(R11415));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11484 (.out1(R11485), .clock(clock), .in1(R11484));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11600 (.out1(R11601), .clock(clock), .in1(R11600));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11661 (.out1(R11662), .clock(clock), .in1(off_3651));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11717 (.out1(R11718), .clock(clock), .in1(_1346));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op1392 (.out1(_1347), .in1(R11718), .in2(1 'd 1));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op1393 (.out1(ifout1393), .in1(_1347), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1461 (.out1(_1415), .in1(R11601));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1454 (.out1(_1408), .in1(R11601));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1443 (.out1(_1397), .in1(R11601));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1423 (.out1(_1377), .in1(R11601));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1462 (.out1(_1416), .in1(_1415), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1455 (.out1(_1409), .in1(_1408), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1444 (.out1(_1398), .in1(_1397), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1424 (.out1(_1378), .in1(_1377), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3877 (.out1(R3878), .clock(clock), .in1(R3877));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4133 (.out1(R4134), .clock(clock), .in1(R4133));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4388 (.out1(R4389), .clock(clock), .in1(R4388));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4633 (.out1(R4634), .clock(clock), .in1(R4633));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4873 (.out1(R4874), .clock(clock), .in1(R4873));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5160 (.out1(R5161), .clock(clock), .in1(R5160));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5392 (.out1(R5393), .clock(clock), .in1(R5392));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5619 (.out1(R5620), .clock(clock), .in1(R5619));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5893 (.out1(R5894), .clock(clock), .in1(R5893));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6111 (.out1(R6112), .clock(clock), .in1(R6111));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6324 (.out1(R6325), .clock(clock), .in1(R6324));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6585 (.out1(R6586), .clock(clock), .in1(R6585));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6790 (.out1(R6791), .clock(clock), .in1(R6790));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6990 (.out1(R6991), .clock(clock), .in1(R6990));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7237 (.out1(R7238), .clock(clock), .in1(R7237));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7429 (.out1(R7430), .clock(clock), .in1(R7429));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7616 (.out1(R7617), .clock(clock), .in1(R7616));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7850 (.out1(R7851), .clock(clock), .in1(R7850));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8029 (.out1(R8030), .clock(clock), .in1(R8029));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8203 (.out1(R8204), .clock(clock), .in1(R8203));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8424 (.out1(R8425), .clock(clock), .in1(R8424));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8590 (.out1(R8591), .clock(clock), .in1(R8590));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8751 (.out1(R8752), .clock(clock), .in1(R8751));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8959 (.out1(R8960), .clock(clock), .in1(R8959));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9112 (.out1(R9113), .clock(clock), .in1(R9112));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9260 (.out1(R9261), .clock(clock), .in1(R9260));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9455 (.out1(R9456), .clock(clock), .in1(R9455));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9595 (.out1(R9596), .clock(clock), .in1(R9595));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9730 (.out1(R9731), .clock(clock), .in1(R9730));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9912 (.out1(R9913), .clock(clock), .in1(R9912));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10039 (.out1(R10040), .clock(clock), .in1(R10039));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10161 (.out1(R10162), .clock(clock), .in1(R10161));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10330 (.out1(R10331), .clock(clock), .in1(R10330));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10443 (.out1(R10444), .clock(clock), .in1(R10443));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10551 (.out1(R10552), .clock(clock), .in1(R10551));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10707 (.out1(R10708), .clock(clock), .in1(R10707));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10807 (.out1(R10808), .clock(clock), .in1(R10807));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10902 (.out1(R10903), .clock(clock), .in1(R10902));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11044 (.out1(R11045), .clock(clock), .in1(R11044));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11131 (.out1(R11132), .clock(clock), .in1(R11131));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11213 (.out1(R11214), .clock(clock), .in1(R11213));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11342 (.out1(R11343), .clock(clock), .in1(R11342));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11416 (.out1(R11417), .clock(clock), .in1(R11416));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11485 (.out1(R11486), .clock(clock), .in1(R11485));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11601 (.out1(R11602), .clock(clock), .in1(R11601));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11662 (.out1(R11663), .clock(clock), .in1(R11662));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11718 (.out1(R11719), .clock(clock), .in1(ifout1393));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11781 (.out1(R11782), .clock(clock), .in1(_1416));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11782 (.out1(R11783), .clock(clock), .in1(_1409));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11783 (.out1(R11784), .clock(clock), .in1(_1398));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11784 (.out1(R11785), .clock(clock), .in1(_1378));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1436 (.out1(_1390), .in1(R11602));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1416 (.out1(_1370), .in1(R11602));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1405 (.out1(_1359), .in1(R11602));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1398 (.out1(_1352), .in1(R11602));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1465 (.out1(_1419), .in1(2 'd 2), .in2(R11663));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1437 (.out1(_1391), .in1(_1390), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1417 (.out1(_1371), .in1(_1370), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1406 (.out1(_1360), .in1(_1359), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1399 (.out1(_1353), .in1(_1352), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1463 (.out1(_1417), .in1(vec100_3652_D), .in2(R11782));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1456 (.out1(_1410), .in1(vec100_3652_D), .in2(R11783));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1445 (.out1(_1399), .in1(vec100_3652_D), .in2(R11784));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1425 (.out1(_1379), .in1(vec100_3652_D), .in2(R11785));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3878 (.out1(R3879), .clock(clock), .in1(R3878));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4134 (.out1(R4135), .clock(clock), .in1(R4134));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4389 (.out1(R4390), .clock(clock), .in1(R4389));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4634 (.out1(R4635), .clock(clock), .in1(R4634));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4874 (.out1(R4875), .clock(clock), .in1(R4874));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5161 (.out1(R5162), .clock(clock), .in1(R5161));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5393 (.out1(R5394), .clock(clock), .in1(R5393));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5620 (.out1(R5621), .clock(clock), .in1(R5620));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5894 (.out1(R5895), .clock(clock), .in1(R5894));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6112 (.out1(R6113), .clock(clock), .in1(R6112));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6325 (.out1(R6326), .clock(clock), .in1(R6325));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6586 (.out1(R6587), .clock(clock), .in1(R6586));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6791 (.out1(R6792), .clock(clock), .in1(R6791));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6991 (.out1(R6992), .clock(clock), .in1(R6991));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7238 (.out1(R7239), .clock(clock), .in1(R7238));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7430 (.out1(R7431), .clock(clock), .in1(R7430));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7617 (.out1(R7618), .clock(clock), .in1(R7617));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7851 (.out1(R7852), .clock(clock), .in1(R7851));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8030 (.out1(R8031), .clock(clock), .in1(R8030));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8204 (.out1(R8205), .clock(clock), .in1(R8204));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8425 (.out1(R8426), .clock(clock), .in1(R8425));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8591 (.out1(R8592), .clock(clock), .in1(R8591));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8752 (.out1(R8753), .clock(clock), .in1(R8752));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8960 (.out1(R8961), .clock(clock), .in1(R8960));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9113 (.out1(R9114), .clock(clock), .in1(R9113));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9261 (.out1(R9262), .clock(clock), .in1(R9261));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9456 (.out1(R9457), .clock(clock), .in1(R9456));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9596 (.out1(R9597), .clock(clock), .in1(R9596));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9731 (.out1(R9732), .clock(clock), .in1(R9731));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9913 (.out1(R9914), .clock(clock), .in1(R9913));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10040 (.out1(R10041), .clock(clock), .in1(R10040));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10162 (.out1(R10163), .clock(clock), .in1(R10162));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10331 (.out1(R10332), .clock(clock), .in1(R10331));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10444 (.out1(R10445), .clock(clock), .in1(R10444));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10552 (.out1(R10553), .clock(clock), .in1(R10552));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10708 (.out1(R10709), .clock(clock), .in1(R10708));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10808 (.out1(R10809), .clock(clock), .in1(R10808));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10903 (.out1(R10904), .clock(clock), .in1(R10903));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11045 (.out1(R11046), .clock(clock), .in1(R11045));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11132 (.out1(R11133), .clock(clock), .in1(R11132));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11214 (.out1(R11215), .clock(clock), .in1(R11214));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11343 (.out1(R11344), .clock(clock), .in1(R11343));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11417 (.out1(R11418), .clock(clock), .in1(R11417));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11486 (.out1(R11487), .clock(clock), .in1(R11486));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11602 (.out1(R11603), .clock(clock), .in1(R11602));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11663 (.out1(R11664), .clock(clock), .in1(R11663));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11719 (.out1(R11720), .clock(clock), .in1(R11719));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11785 (.out1(R11786), .clock(clock), .in1(_1419));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11786 (.out1(R11787), .clock(clock), .in1(_1391));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11787 (.out1(R11788), .clock(clock), .in1(_1371));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11788 (.out1(R11789), .clock(clock), .in1(_1360));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11789 (.out1(R11790), .clock(clock), .in1(_1353));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11790 (.out1(R11791), .clock(clock), .in1(_1417));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11791 (.out1(R11792), .clock(clock), .in1(_1410));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11792 (.out1(R11793), .clock(clock), .in1(_1399));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11793 (.out1(R11794), .clock(clock), .in1(_1379));
  SRAM op1464 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1418),.ADR(R11791));
  SRAM op1457 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1411),.ADR(R11792));
  SRAM op1446 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1400),.ADR(R11793));
  SRAM op1426 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1380),.ADR(R11794));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1458 (.out1(_1412), .in1(2 'd 2), .in2(R11664));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1447 (.out1(_1401), .in1(2 'd 2), .in2(R11664));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1440 (.out1(_1394), .in1(2 'd 2), .in2(R11664));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1427 (.out1(_1381), .in1(2 'd 2), .in2(R11664));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1420 (.out1(_1374), .in1(2 'd 2), .in2(R11664));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1409 (.out1(_1363), .in1(2 'd 2), .in2(R11664));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1438 (.out1(_1392), .in1(vec100_3652_D), .in2(R11787));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1418 (.out1(_1372), .in1(vec100_3652_D), .in2(R11788));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1407 (.out1(_1361), .in1(vec100_3652_D), .in2(R11789));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1400 (.out1(_1354), .in1(vec100_3652_D), .in2(R11790));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1466 (.out1(_1420), .in1(R11786), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3879 (.out1(R3880), .clock(clock), .in1(R3879));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4135 (.out1(R4136), .clock(clock), .in1(R4135));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4390 (.out1(R4391), .clock(clock), .in1(R4390));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4635 (.out1(R4636), .clock(clock), .in1(R4635));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4875 (.out1(R4876), .clock(clock), .in1(R4875));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5162 (.out1(R5163), .clock(clock), .in1(R5162));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5394 (.out1(R5395), .clock(clock), .in1(R5394));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5621 (.out1(R5622), .clock(clock), .in1(R5621));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5895 (.out1(R5896), .clock(clock), .in1(R5895));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6113 (.out1(R6114), .clock(clock), .in1(R6113));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6326 (.out1(R6327), .clock(clock), .in1(R6326));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6587 (.out1(R6588), .clock(clock), .in1(R6587));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6792 (.out1(R6793), .clock(clock), .in1(R6792));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6992 (.out1(R6993), .clock(clock), .in1(R6992));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7239 (.out1(R7240), .clock(clock), .in1(R7239));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7431 (.out1(R7432), .clock(clock), .in1(R7431));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7618 (.out1(R7619), .clock(clock), .in1(R7618));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7852 (.out1(R7853), .clock(clock), .in1(R7852));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8031 (.out1(R8032), .clock(clock), .in1(R8031));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8205 (.out1(R8206), .clock(clock), .in1(R8205));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8426 (.out1(R8427), .clock(clock), .in1(R8426));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8592 (.out1(R8593), .clock(clock), .in1(R8592));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8753 (.out1(R8754), .clock(clock), .in1(R8753));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8961 (.out1(R8962), .clock(clock), .in1(R8961));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9114 (.out1(R9115), .clock(clock), .in1(R9114));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9262 (.out1(R9263), .clock(clock), .in1(R9262));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9457 (.out1(R9458), .clock(clock), .in1(R9457));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9597 (.out1(R9598), .clock(clock), .in1(R9597));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9732 (.out1(R9733), .clock(clock), .in1(R9732));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9914 (.out1(R9915), .clock(clock), .in1(R9914));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10041 (.out1(R10042), .clock(clock), .in1(R10041));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10163 (.out1(R10164), .clock(clock), .in1(R10163));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10332 (.out1(R10333), .clock(clock), .in1(R10332));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10445 (.out1(R10446), .clock(clock), .in1(R10445));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10553 (.out1(R10554), .clock(clock), .in1(R10553));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10709 (.out1(R10710), .clock(clock), .in1(R10709));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10809 (.out1(R10810), .clock(clock), .in1(R10809));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10904 (.out1(R10905), .clock(clock), .in1(R10904));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11046 (.out1(R11047), .clock(clock), .in1(R11046));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11133 (.out1(R11134), .clock(clock), .in1(R11133));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11215 (.out1(R11216), .clock(clock), .in1(R11215));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11344 (.out1(R11345), .clock(clock), .in1(R11344));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11418 (.out1(R11419), .clock(clock), .in1(R11418));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11487 (.out1(R11488), .clock(clock), .in1(R11487));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11603 (.out1(R11604), .clock(clock), .in1(R11603));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11664 (.out1(R11665), .clock(clock), .in1(R11664));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11720 (.out1(R11721), .clock(clock), .in1(R11720));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11794 (.out1(R11795), .clock(clock), .in1(_1418));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11795 (.out1(R11796), .clock(clock), .in1(_1411));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11796 (.out1(R11797), .clock(clock), .in1(_1400));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11797 (.out1(R11798), .clock(clock), .in1(_1380));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11798 (.out1(R11799), .clock(clock), .in1(_1412));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11799 (.out1(R11800), .clock(clock), .in1(_1401));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11800 (.out1(R11801), .clock(clock), .in1(_1394));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11801 (.out1(R11802), .clock(clock), .in1(_1381));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11802 (.out1(R11803), .clock(clock), .in1(_1374));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11803 (.out1(R11804), .clock(clock), .in1(_1363));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11804 (.out1(R11805), .clock(clock), .in1(_1392));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11805 (.out1(R11806), .clock(clock), .in1(_1372));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11806 (.out1(R11807), .clock(clock), .in1(_1361));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11807 (.out1(R11808), .clock(clock), .in1(_1354));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11808 (.out1(R11809), .clock(clock), .in1(_1420));
  SRAM op1439 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1393),.ADR(R11805));
  SRAM op1419 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1373),.ADR(R11806));
  SRAM op1408 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1362),.ADR(R11807));
  SRAM op1401 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1355),.ADR(R11808));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1467 (.out1(_1421), .in1(R11795), .in2(R11809));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1468 (.out1(_1422), .in1(_1421), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1459 (.out1(_1413), .in1(R11799), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1448 (.out1(_1402), .in1(R11800), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1428 (.out1(_1382), .in1(R11802), .in2(64 'd 18446744073709551615));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1402 (.out1(_1356), .in1(2 'd 2), .in2(R11665));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1469 (.out1(_1423), .in1(_1422), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1460 (.out1(_1414), .in1(R11796), .in2(_1413));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1449 (.out1(_1403), .in1(R11797), .in2(_1402));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1429 (.out1(_1383), .in1(R11798), .in2(_1382));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1470 (.out1(_1424), .in1(_1414), .in2(_1423));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1450 (.out1(_1404), .in1(_1403), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1441 (.out1(_1395), .in1(R11801), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1430 (.out1(_1384), .in1(_1383), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1421 (.out1(_1375), .in1(R11803), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1410 (.out1(_1364), .in1(R11804), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3880 (.out1(R3881), .clock(clock), .in1(R3880));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4136 (.out1(R4137), .clock(clock), .in1(R4136));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4391 (.out1(R4392), .clock(clock), .in1(R4391));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4636 (.out1(R4637), .clock(clock), .in1(R4636));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4876 (.out1(R4877), .clock(clock), .in1(R4876));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5163 (.out1(R5164), .clock(clock), .in1(R5163));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5395 (.out1(R5396), .clock(clock), .in1(R5395));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5622 (.out1(R5623), .clock(clock), .in1(R5622));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5896 (.out1(R5897), .clock(clock), .in1(R5896));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6114 (.out1(R6115), .clock(clock), .in1(R6114));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6327 (.out1(R6328), .clock(clock), .in1(R6327));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6588 (.out1(R6589), .clock(clock), .in1(R6588));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6793 (.out1(R6794), .clock(clock), .in1(R6793));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6993 (.out1(R6994), .clock(clock), .in1(R6993));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7240 (.out1(R7241), .clock(clock), .in1(R7240));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7432 (.out1(R7433), .clock(clock), .in1(R7432));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7619 (.out1(R7620), .clock(clock), .in1(R7619));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7853 (.out1(R7854), .clock(clock), .in1(R7853));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8032 (.out1(R8033), .clock(clock), .in1(R8032));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8206 (.out1(R8207), .clock(clock), .in1(R8206));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8427 (.out1(R8428), .clock(clock), .in1(R8427));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8593 (.out1(R8594), .clock(clock), .in1(R8593));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8754 (.out1(R8755), .clock(clock), .in1(R8754));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8962 (.out1(R8963), .clock(clock), .in1(R8962));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9115 (.out1(R9116), .clock(clock), .in1(R9115));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9263 (.out1(R9264), .clock(clock), .in1(R9263));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9458 (.out1(R9459), .clock(clock), .in1(R9458));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9598 (.out1(R9599), .clock(clock), .in1(R9598));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9733 (.out1(R9734), .clock(clock), .in1(R9733));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9915 (.out1(R9916), .clock(clock), .in1(R9915));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10042 (.out1(R10043), .clock(clock), .in1(R10042));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10164 (.out1(R10165), .clock(clock), .in1(R10164));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10333 (.out1(R10334), .clock(clock), .in1(R10333));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10446 (.out1(R10447), .clock(clock), .in1(R10446));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10554 (.out1(R10555), .clock(clock), .in1(R10554));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10710 (.out1(R10711), .clock(clock), .in1(R10710));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10810 (.out1(R10811), .clock(clock), .in1(R10810));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10905 (.out1(R10906), .clock(clock), .in1(R10905));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11047 (.out1(R11048), .clock(clock), .in1(R11047));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11134 (.out1(R11135), .clock(clock), .in1(R11134));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11216 (.out1(R11217), .clock(clock), .in1(R11216));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11345 (.out1(R11346), .clock(clock), .in1(R11345));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11419 (.out1(R11420), .clock(clock), .in1(R11419));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11488 (.out1(R11489), .clock(clock), .in1(R11488));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11604 (.out1(R11605), .clock(clock), .in1(R11604));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11665 (.out1(R11666), .clock(clock), .in1(R11665));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11721 (.out1(R11722), .clock(clock), .in1(R11721));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11809 (.out1(R11810), .clock(clock), .in1(_1393));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11810 (.out1(R11811), .clock(clock), .in1(_1373));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11811 (.out1(R11812), .clock(clock), .in1(_1362));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11812 (.out1(R11813), .clock(clock), .in1(_1355));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11813 (.out1(R11814), .clock(clock), .in1(_1356));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11814 (.out1(R11815), .clock(clock), .in1(_1424));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11815 (.out1(R11816), .clock(clock), .in1(_1404));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11816 (.out1(R11817), .clock(clock), .in1(_1395));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11817 (.out1(R11818), .clock(clock), .in1(_1384));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11818 (.out1(R11819), .clock(clock), .in1(_1375));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11819 (.out1(R11820), .clock(clock), .in1(_1364));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1451 (.out1(_1405), .in1(R11816), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1442 (.out1(_1396), .in1(R11810), .in2(R11817));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1411 (.out1(_1365), .in1(R11812), .in2(R11820));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1471 (.out1(_1425), .in1(R11815), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1452 (.out1(_1406), .in1(_1396), .in2(_1405));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1431 (.out1(_1385), .in1(R11818), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1422 (.out1(_1376), .in1(R11811), .in2(R11819));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1412 (.out1(_1366), .in1(_1365), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1403 (.out1(_1357), .in1(R11814), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1432 (.out1(_1386), .in1(_1376), .in2(_1385));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1472 (.out1(_1426), .in1(_1425), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1453 (.out1(_1407), .in1(_1406), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1413 (.out1(_1367), .in1(_1366), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1404 (.out1(_1358), .in1(R11813), .in2(_1357));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1473 (.out1(_1427), .in1(_1407), .in2(_1426));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1433 (.out1(_1387), .in1(_1386), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1414 (.out1(_1368), .in1(_1358), .in2(_1367));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3881 (.out1(R3882), .clock(clock), .in1(R3881));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4137 (.out1(R4138), .clock(clock), .in1(R4137));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4392 (.out1(R4393), .clock(clock), .in1(R4392));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4637 (.out1(R4638), .clock(clock), .in1(R4637));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4877 (.out1(R4878), .clock(clock), .in1(R4877));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5164 (.out1(R5165), .clock(clock), .in1(R5164));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5396 (.out1(R5397), .clock(clock), .in1(R5396));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5623 (.out1(R5624), .clock(clock), .in1(R5623));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5897 (.out1(R5898), .clock(clock), .in1(R5897));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6115 (.out1(R6116), .clock(clock), .in1(R6115));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6328 (.out1(R6329), .clock(clock), .in1(R6328));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6589 (.out1(R6590), .clock(clock), .in1(R6589));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6794 (.out1(R6795), .clock(clock), .in1(R6794));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6994 (.out1(R6995), .clock(clock), .in1(R6994));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7241 (.out1(R7242), .clock(clock), .in1(R7241));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7433 (.out1(R7434), .clock(clock), .in1(R7433));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7620 (.out1(R7621), .clock(clock), .in1(R7620));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7854 (.out1(R7855), .clock(clock), .in1(R7854));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8033 (.out1(R8034), .clock(clock), .in1(R8033));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8207 (.out1(R8208), .clock(clock), .in1(R8207));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8428 (.out1(R8429), .clock(clock), .in1(R8428));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8594 (.out1(R8595), .clock(clock), .in1(R8594));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8755 (.out1(R8756), .clock(clock), .in1(R8755));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8963 (.out1(R8964), .clock(clock), .in1(R8963));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9116 (.out1(R9117), .clock(clock), .in1(R9116));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9264 (.out1(R9265), .clock(clock), .in1(R9264));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9459 (.out1(R9460), .clock(clock), .in1(R9459));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9599 (.out1(R9600), .clock(clock), .in1(R9599));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9734 (.out1(R9735), .clock(clock), .in1(R9734));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9916 (.out1(R9917), .clock(clock), .in1(R9916));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10043 (.out1(R10044), .clock(clock), .in1(R10043));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10165 (.out1(R10166), .clock(clock), .in1(R10165));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10334 (.out1(R10335), .clock(clock), .in1(R10334));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10447 (.out1(R10448), .clock(clock), .in1(R10447));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10555 (.out1(R10556), .clock(clock), .in1(R10555));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10711 (.out1(R10712), .clock(clock), .in1(R10711));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10811 (.out1(R10812), .clock(clock), .in1(R10811));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10906 (.out1(R10907), .clock(clock), .in1(R10906));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11048 (.out1(R11049), .clock(clock), .in1(R11048));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11135 (.out1(R11136), .clock(clock), .in1(R11135));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11217 (.out1(R11218), .clock(clock), .in1(R11217));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11346 (.out1(R11347), .clock(clock), .in1(R11346));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11420 (.out1(R11421), .clock(clock), .in1(R11420));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11489 (.out1(R11490), .clock(clock), .in1(R11489));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11605 (.out1(R11606), .clock(clock), .in1(R11605));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11666 (.out1(R11667), .clock(clock), .in1(R11666));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11722 (.out1(R11723), .clock(clock), .in1(R11722));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11820 (.out1(R11821), .clock(clock), .in1(_1427));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11821 (.out1(R11822), .clock(clock), .in1(_1387));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11822 (.out1(R11823), .clock(clock), .in1(_1368));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1394 (.out1(_1348), .in1(R11606));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1434 (.out1(_1388), .in1(R11822), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1415 (.out1(_1369), .in1(R11823), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op1474 (.out1(_1428), .in1(R11821), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1435 (.out1(_1389), .in1(_1369), .in2(_1388));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1395 (.out1(_1349), .in1(_1348), .in2(2 'd 2));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1475 (.out1(_1429), .in1(_1389), .in2(_1428));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op1476 (.out1(_1430), .in1(_1429), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3882 (.out1(R3883), .clock(clock), .in1(R3882));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4138 (.out1(R4139), .clock(clock), .in1(R4138));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4393 (.out1(R4394), .clock(clock), .in1(R4393));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4638 (.out1(R4639), .clock(clock), .in1(R4638));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4878 (.out1(R4879), .clock(clock), .in1(R4878));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5165 (.out1(R5166), .clock(clock), .in1(R5165));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5397 (.out1(R5398), .clock(clock), .in1(R5397));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5624 (.out1(R5625), .clock(clock), .in1(R5624));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5898 (.out1(R5899), .clock(clock), .in1(R5898));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6116 (.out1(R6117), .clock(clock), .in1(R6116));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6329 (.out1(R6330), .clock(clock), .in1(R6329));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6590 (.out1(R6591), .clock(clock), .in1(R6590));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6795 (.out1(R6796), .clock(clock), .in1(R6795));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6995 (.out1(R6996), .clock(clock), .in1(R6995));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7242 (.out1(R7243), .clock(clock), .in1(R7242));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7434 (.out1(R7435), .clock(clock), .in1(R7434));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7621 (.out1(R7622), .clock(clock), .in1(R7621));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7855 (.out1(R7856), .clock(clock), .in1(R7855));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8034 (.out1(R8035), .clock(clock), .in1(R8034));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8208 (.out1(R8209), .clock(clock), .in1(R8208));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8429 (.out1(R8430), .clock(clock), .in1(R8429));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8595 (.out1(R8596), .clock(clock), .in1(R8595));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8756 (.out1(R8757), .clock(clock), .in1(R8756));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8964 (.out1(R8965), .clock(clock), .in1(R8964));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9117 (.out1(R9118), .clock(clock), .in1(R9117));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9265 (.out1(R9266), .clock(clock), .in1(R9265));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9460 (.out1(R9461), .clock(clock), .in1(R9460));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9600 (.out1(R9601), .clock(clock), .in1(R9600));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9735 (.out1(R9736), .clock(clock), .in1(R9735));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9917 (.out1(R9918), .clock(clock), .in1(R9917));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10044 (.out1(R10045), .clock(clock), .in1(R10044));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10166 (.out1(R10167), .clock(clock), .in1(R10166));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10335 (.out1(R10336), .clock(clock), .in1(R10335));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10448 (.out1(R10449), .clock(clock), .in1(R10448));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10556 (.out1(R10557), .clock(clock), .in1(R10556));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10712 (.out1(R10713), .clock(clock), .in1(R10712));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10812 (.out1(R10813), .clock(clock), .in1(R10812));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10907 (.out1(R10908), .clock(clock), .in1(R10907));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11049 (.out1(R11050), .clock(clock), .in1(R11049));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11136 (.out1(R11137), .clock(clock), .in1(R11136));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11218 (.out1(R11219), .clock(clock), .in1(R11218));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11347 (.out1(R11348), .clock(clock), .in1(R11347));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11421 (.out1(R11422), .clock(clock), .in1(R11421));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11490 (.out1(R11491), .clock(clock), .in1(R11490));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11606 (.out1(R11607), .clock(clock), .in1(R11606));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11667 (.out1(R11668), .clock(clock), .in1(R11667));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11723 (.out1(R11724), .clock(clock), .in1(R11723));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11823 (.out1(R11824), .clock(clock), .in1(_1349));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11824 (.out1(R11825), .clock(clock), .in1(_1430));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op1477 (.out1(_1431), .in1(R11825), .in2(57 'd 72340172838076673));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1396 (.out1(_1350), .in1(base0_100_3657_D), .in2(R11824));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3883 (.out1(R3884), .clock(clock), .in1(R3883));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4139 (.out1(R4140), .clock(clock), .in1(R4139));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4394 (.out1(R4395), .clock(clock), .in1(R4394));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4639 (.out1(R4640), .clock(clock), .in1(R4639));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4879 (.out1(R4880), .clock(clock), .in1(R4879));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5166 (.out1(R5167), .clock(clock), .in1(R5166));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5398 (.out1(R5399), .clock(clock), .in1(R5398));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5625 (.out1(R5626), .clock(clock), .in1(R5625));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5899 (.out1(R5900), .clock(clock), .in1(R5899));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6117 (.out1(R6118), .clock(clock), .in1(R6117));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6330 (.out1(R6331), .clock(clock), .in1(R6330));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6591 (.out1(R6592), .clock(clock), .in1(R6591));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6796 (.out1(R6797), .clock(clock), .in1(R6796));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6996 (.out1(R6997), .clock(clock), .in1(R6996));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7243 (.out1(R7244), .clock(clock), .in1(R7243));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7435 (.out1(R7436), .clock(clock), .in1(R7435));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7622 (.out1(R7623), .clock(clock), .in1(R7622));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7856 (.out1(R7857), .clock(clock), .in1(R7856));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8035 (.out1(R8036), .clock(clock), .in1(R8035));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8209 (.out1(R8210), .clock(clock), .in1(R8209));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8430 (.out1(R8431), .clock(clock), .in1(R8430));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8596 (.out1(R8597), .clock(clock), .in1(R8596));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8757 (.out1(R8758), .clock(clock), .in1(R8757));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8965 (.out1(R8966), .clock(clock), .in1(R8965));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9118 (.out1(R9119), .clock(clock), .in1(R9118));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9266 (.out1(R9267), .clock(clock), .in1(R9266));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9461 (.out1(R9462), .clock(clock), .in1(R9461));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9601 (.out1(R9602), .clock(clock), .in1(R9601));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9736 (.out1(R9737), .clock(clock), .in1(R9736));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9918 (.out1(R9919), .clock(clock), .in1(R9918));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10045 (.out1(R10046), .clock(clock), .in1(R10045));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10167 (.out1(R10168), .clock(clock), .in1(R10167));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10336 (.out1(R10337), .clock(clock), .in1(R10336));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10449 (.out1(R10450), .clock(clock), .in1(R10449));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10557 (.out1(R10558), .clock(clock), .in1(R10557));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10713 (.out1(R10714), .clock(clock), .in1(R10713));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10813 (.out1(R10814), .clock(clock), .in1(R10813));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10908 (.out1(R10909), .clock(clock), .in1(R10908));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11050 (.out1(R11051), .clock(clock), .in1(R11050));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11137 (.out1(R11138), .clock(clock), .in1(R11137));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11219 (.out1(R11220), .clock(clock), .in1(R11219));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11348 (.out1(R11349), .clock(clock), .in1(R11348));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11422 (.out1(R11423), .clock(clock), .in1(R11422));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11491 (.out1(R11492), .clock(clock), .in1(R11491));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11607 (.out1(R11608), .clock(clock), .in1(R11607));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11668 (.out1(R11669), .clock(clock), .in1(R11668));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11724 (.out1(R11725), .clock(clock), .in1(R11724));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11825 (.out1(R11826), .clock(clock), .in1(_1431));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11826 (.out1(R11827), .clock(clock), .in1(_1350));
  SRAM op1397 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1351),.ADR(R11827));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op1478 (.out1(_1432), .in1(R11826), .in2(6 'd 56));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3884 (.out1(R3885), .clock(clock), .in1(R3884));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4140 (.out1(R4141), .clock(clock), .in1(R4140));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4395 (.out1(R4396), .clock(clock), .in1(R4395));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4640 (.out1(R4641), .clock(clock), .in1(R4640));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4880 (.out1(R4881), .clock(clock), .in1(R4880));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5167 (.out1(R5168), .clock(clock), .in1(R5167));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5399 (.out1(R5400), .clock(clock), .in1(R5399));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5626 (.out1(R5627), .clock(clock), .in1(R5626));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5900 (.out1(R5901), .clock(clock), .in1(R5900));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6118 (.out1(R6119), .clock(clock), .in1(R6118));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6331 (.out1(R6332), .clock(clock), .in1(R6331));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6592 (.out1(R6593), .clock(clock), .in1(R6592));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6797 (.out1(R6798), .clock(clock), .in1(R6797));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6997 (.out1(R6998), .clock(clock), .in1(R6997));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7244 (.out1(R7245), .clock(clock), .in1(R7244));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7436 (.out1(R7437), .clock(clock), .in1(R7436));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7623 (.out1(R7624), .clock(clock), .in1(R7623));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7857 (.out1(R7858), .clock(clock), .in1(R7857));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8036 (.out1(R8037), .clock(clock), .in1(R8036));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8210 (.out1(R8211), .clock(clock), .in1(R8210));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8431 (.out1(R8432), .clock(clock), .in1(R8431));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8597 (.out1(R8598), .clock(clock), .in1(R8597));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8758 (.out1(R8759), .clock(clock), .in1(R8758));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8966 (.out1(R8967), .clock(clock), .in1(R8966));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9119 (.out1(R9120), .clock(clock), .in1(R9119));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9267 (.out1(R9268), .clock(clock), .in1(R9267));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9462 (.out1(R9463), .clock(clock), .in1(R9462));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9602 (.out1(R9603), .clock(clock), .in1(R9602));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9737 (.out1(R9738), .clock(clock), .in1(R9737));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9919 (.out1(R9920), .clock(clock), .in1(R9919));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10046 (.out1(R10047), .clock(clock), .in1(R10046));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10168 (.out1(R10169), .clock(clock), .in1(R10168));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10337 (.out1(R10338), .clock(clock), .in1(R10337));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10450 (.out1(R10451), .clock(clock), .in1(R10450));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10558 (.out1(R10559), .clock(clock), .in1(R10558));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10714 (.out1(R10715), .clock(clock), .in1(R10714));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10814 (.out1(R10815), .clock(clock), .in1(R10814));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10909 (.out1(R10910), .clock(clock), .in1(R10909));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11051 (.out1(R11052), .clock(clock), .in1(R11051));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11138 (.out1(R11139), .clock(clock), .in1(R11138));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11220 (.out1(R11221), .clock(clock), .in1(R11220));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11349 (.out1(R11350), .clock(clock), .in1(R11349));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11423 (.out1(R11424), .clock(clock), .in1(R11423));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11492 (.out1(R11493), .clock(clock), .in1(R11492));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11608 (.out1(R11609), .clock(clock), .in1(R11608));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11669 (.out1(R11670), .clock(clock), .in1(R11669));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11725 (.out1(R11726), .clock(clock), .in1(R11725));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11827 (.out1(R11828), .clock(clock), .in1(_1351));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11828 (.out1(R11829), .clock(clock), .in1(_1432));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1479 (.out1(_1433), .in1(R11829));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1480 (.out1(_1434), .in1(R11828), .in2(_1433));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1481 (.out1(idx_3658), .in1(_1434), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3885 (.out1(R3886), .clock(clock), .in1(R3885));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4141 (.out1(R4142), .clock(clock), .in1(R4141));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4396 (.out1(R4397), .clock(clock), .in1(R4396));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4641 (.out1(R4642), .clock(clock), .in1(R4641));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4881 (.out1(R4882), .clock(clock), .in1(R4881));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5168 (.out1(R5169), .clock(clock), .in1(R5168));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5400 (.out1(R5401), .clock(clock), .in1(R5400));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5627 (.out1(R5628), .clock(clock), .in1(R5627));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5901 (.out1(R5902), .clock(clock), .in1(R5901));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6119 (.out1(R6120), .clock(clock), .in1(R6119));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6332 (.out1(R6333), .clock(clock), .in1(R6332));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6593 (.out1(R6594), .clock(clock), .in1(R6593));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6798 (.out1(R6799), .clock(clock), .in1(R6798));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6998 (.out1(R6999), .clock(clock), .in1(R6998));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7245 (.out1(R7246), .clock(clock), .in1(R7245));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7437 (.out1(R7438), .clock(clock), .in1(R7437));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7624 (.out1(R7625), .clock(clock), .in1(R7624));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7858 (.out1(R7859), .clock(clock), .in1(R7858));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8037 (.out1(R8038), .clock(clock), .in1(R8037));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8211 (.out1(R8212), .clock(clock), .in1(R8211));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8432 (.out1(R8433), .clock(clock), .in1(R8432));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8598 (.out1(R8599), .clock(clock), .in1(R8598));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8759 (.out1(R8760), .clock(clock), .in1(R8759));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8967 (.out1(R8968), .clock(clock), .in1(R8967));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9120 (.out1(R9121), .clock(clock), .in1(R9120));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9268 (.out1(R9269), .clock(clock), .in1(R9268));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9463 (.out1(R9464), .clock(clock), .in1(R9463));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9603 (.out1(R9604), .clock(clock), .in1(R9603));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9738 (.out1(R9739), .clock(clock), .in1(R9738));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9920 (.out1(R9921), .clock(clock), .in1(R9920));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10047 (.out1(R10048), .clock(clock), .in1(R10047));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10169 (.out1(R10170), .clock(clock), .in1(R10169));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10338 (.out1(R10339), .clock(clock), .in1(R10338));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10451 (.out1(R10452), .clock(clock), .in1(R10451));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10559 (.out1(R10560), .clock(clock), .in1(R10559));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10715 (.out1(R10716), .clock(clock), .in1(R10715));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10815 (.out1(R10816), .clock(clock), .in1(R10815));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10910 (.out1(R10911), .clock(clock), .in1(R10910));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11052 (.out1(R11053), .clock(clock), .in1(R11052));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11139 (.out1(R11140), .clock(clock), .in1(R11139));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11221 (.out1(R11222), .clock(clock), .in1(R11221));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11350 (.out1(R11351), .clock(clock), .in1(R11350));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11424 (.out1(R11425), .clock(clock), .in1(R11424));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11493 (.out1(R11494), .clock(clock), .in1(R11493));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11609 (.out1(R11610), .clock(clock), .in1(R11609));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11670 (.out1(R11671), .clock(clock), .in1(R11670));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11726 (.out1(R11727), .clock(clock), .in1(R11726));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11829 (.out1(R11830), .clock(clock), .in1(idx_3658));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1485 (.out1(_1437), .in1(R11830));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1486 (.out1(_1438), .in1(_1437), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3886 (.out1(R3887), .clock(clock), .in1(R3886));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4142 (.out1(R4143), .clock(clock), .in1(R4142));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4397 (.out1(R4398), .clock(clock), .in1(R4397));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4642 (.out1(R4643), .clock(clock), .in1(R4642));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4882 (.out1(R4883), .clock(clock), .in1(R4882));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5169 (.out1(R5170), .clock(clock), .in1(R5169));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5401 (.out1(R5402), .clock(clock), .in1(R5401));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5628 (.out1(R5629), .clock(clock), .in1(R5628));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5902 (.out1(R5903), .clock(clock), .in1(R5902));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6120 (.out1(R6121), .clock(clock), .in1(R6120));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6333 (.out1(R6334), .clock(clock), .in1(R6333));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6594 (.out1(R6595), .clock(clock), .in1(R6594));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6799 (.out1(R6800), .clock(clock), .in1(R6799));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6999 (.out1(R7000), .clock(clock), .in1(R6999));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7246 (.out1(R7247), .clock(clock), .in1(R7246));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7438 (.out1(R7439), .clock(clock), .in1(R7438));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7625 (.out1(R7626), .clock(clock), .in1(R7625));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7859 (.out1(R7860), .clock(clock), .in1(R7859));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8038 (.out1(R8039), .clock(clock), .in1(R8038));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8212 (.out1(R8213), .clock(clock), .in1(R8212));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8433 (.out1(R8434), .clock(clock), .in1(R8433));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8599 (.out1(R8600), .clock(clock), .in1(R8599));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8760 (.out1(R8761), .clock(clock), .in1(R8760));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8968 (.out1(R8969), .clock(clock), .in1(R8968));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9121 (.out1(R9122), .clock(clock), .in1(R9121));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9269 (.out1(R9270), .clock(clock), .in1(R9269));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9464 (.out1(R9465), .clock(clock), .in1(R9464));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9604 (.out1(R9605), .clock(clock), .in1(R9604));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9739 (.out1(R9740), .clock(clock), .in1(R9739));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9921 (.out1(R9922), .clock(clock), .in1(R9921));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10048 (.out1(R10049), .clock(clock), .in1(R10048));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10170 (.out1(R10171), .clock(clock), .in1(R10170));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10339 (.out1(R10340), .clock(clock), .in1(R10339));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10452 (.out1(R10453), .clock(clock), .in1(R10452));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10560 (.out1(R10561), .clock(clock), .in1(R10560));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10716 (.out1(R10717), .clock(clock), .in1(R10716));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10816 (.out1(R10817), .clock(clock), .in1(R10816));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10911 (.out1(R10912), .clock(clock), .in1(R10911));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11053 (.out1(R11054), .clock(clock), .in1(R11053));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11140 (.out1(R11141), .clock(clock), .in1(R11140));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11222 (.out1(R11223), .clock(clock), .in1(R11222));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11351 (.out1(R11352), .clock(clock), .in1(R11351));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11425 (.out1(R11426), .clock(clock), .in1(R11425));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11494 (.out1(R11495), .clock(clock), .in1(R11494));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11610 (.out1(R11611), .clock(clock), .in1(R11610));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11671 (.out1(R11672), .clock(clock), .in1(R11671));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11727 (.out1(R11728), .clock(clock), .in1(R11727));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11830 (.out1(R11831), .clock(clock), .in1(R11830));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11878 (.out1(R11879), .clock(clock), .in1(_1438));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1487 (.out1(_1439), .in1(vec106_3660_D), .in2(R11879));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3887 (.out1(R3888), .clock(clock), .in1(R3887));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4143 (.out1(R4144), .clock(clock), .in1(R4143));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4398 (.out1(R4399), .clock(clock), .in1(R4398));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4643 (.out1(R4644), .clock(clock), .in1(R4643));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4883 (.out1(R4884), .clock(clock), .in1(R4883));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5170 (.out1(R5171), .clock(clock), .in1(R5170));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5402 (.out1(R5403), .clock(clock), .in1(R5402));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5629 (.out1(R5630), .clock(clock), .in1(R5629));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5903 (.out1(R5904), .clock(clock), .in1(R5903));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6121 (.out1(R6122), .clock(clock), .in1(R6121));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6334 (.out1(R6335), .clock(clock), .in1(R6334));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6595 (.out1(R6596), .clock(clock), .in1(R6595));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6800 (.out1(R6801), .clock(clock), .in1(R6800));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7000 (.out1(R7001), .clock(clock), .in1(R7000));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7247 (.out1(R7248), .clock(clock), .in1(R7247));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7439 (.out1(R7440), .clock(clock), .in1(R7439));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7626 (.out1(R7627), .clock(clock), .in1(R7626));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7860 (.out1(R7861), .clock(clock), .in1(R7860));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8039 (.out1(R8040), .clock(clock), .in1(R8039));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8213 (.out1(R8214), .clock(clock), .in1(R8213));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8434 (.out1(R8435), .clock(clock), .in1(R8434));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8600 (.out1(R8601), .clock(clock), .in1(R8600));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8761 (.out1(R8762), .clock(clock), .in1(R8761));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8969 (.out1(R8970), .clock(clock), .in1(R8969));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9122 (.out1(R9123), .clock(clock), .in1(R9122));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9270 (.out1(R9271), .clock(clock), .in1(R9270));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9465 (.out1(R9466), .clock(clock), .in1(R9465));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9605 (.out1(R9606), .clock(clock), .in1(R9605));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9740 (.out1(R9741), .clock(clock), .in1(R9740));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9922 (.out1(R9923), .clock(clock), .in1(R9922));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10049 (.out1(R10050), .clock(clock), .in1(R10049));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10171 (.out1(R10172), .clock(clock), .in1(R10171));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10340 (.out1(R10341), .clock(clock), .in1(R10340));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10453 (.out1(R10454), .clock(clock), .in1(R10453));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10561 (.out1(R10562), .clock(clock), .in1(R10561));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10717 (.out1(R10718), .clock(clock), .in1(R10717));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10817 (.out1(R10818), .clock(clock), .in1(R10817));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10912 (.out1(R10913), .clock(clock), .in1(R10912));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11054 (.out1(R11055), .clock(clock), .in1(R11054));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11141 (.out1(R11142), .clock(clock), .in1(R11141));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11223 (.out1(R11224), .clock(clock), .in1(R11223));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11352 (.out1(R11353), .clock(clock), .in1(R11352));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11426 (.out1(R11427), .clock(clock), .in1(R11426));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11495 (.out1(R11496), .clock(clock), .in1(R11495));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11611 (.out1(R11612), .clock(clock), .in1(R11611));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11672 (.out1(R11673), .clock(clock), .in1(R11672));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11728 (.out1(R11729), .clock(clock), .in1(R11728));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11831 (.out1(R11832), .clock(clock), .in1(R11831));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11879 (.out1(R11880), .clock(clock), .in1(_1439));
  SRAM op1488 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1440),.ADR(R11880));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3888 (.out1(R3889), .clock(clock), .in1(R3888));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4144 (.out1(R4145), .clock(clock), .in1(R4144));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4399 (.out1(R4400), .clock(clock), .in1(R4399));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4644 (.out1(R4645), .clock(clock), .in1(R4644));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4884 (.out1(R4885), .clock(clock), .in1(R4884));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5171 (.out1(R5172), .clock(clock), .in1(R5171));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5403 (.out1(R5404), .clock(clock), .in1(R5403));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5630 (.out1(R5631), .clock(clock), .in1(R5630));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5904 (.out1(R5905), .clock(clock), .in1(R5904));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6122 (.out1(R6123), .clock(clock), .in1(R6122));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6335 (.out1(R6336), .clock(clock), .in1(R6335));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6596 (.out1(R6597), .clock(clock), .in1(R6596));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6801 (.out1(R6802), .clock(clock), .in1(R6801));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7001 (.out1(R7002), .clock(clock), .in1(R7001));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7248 (.out1(R7249), .clock(clock), .in1(R7248));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7440 (.out1(R7441), .clock(clock), .in1(R7440));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7627 (.out1(R7628), .clock(clock), .in1(R7627));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7861 (.out1(R7862), .clock(clock), .in1(R7861));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8040 (.out1(R8041), .clock(clock), .in1(R8040));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8214 (.out1(R8215), .clock(clock), .in1(R8214));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8435 (.out1(R8436), .clock(clock), .in1(R8435));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8601 (.out1(R8602), .clock(clock), .in1(R8601));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8762 (.out1(R8763), .clock(clock), .in1(R8762));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8970 (.out1(R8971), .clock(clock), .in1(R8970));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9123 (.out1(R9124), .clock(clock), .in1(R9123));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9271 (.out1(R9272), .clock(clock), .in1(R9271));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9466 (.out1(R9467), .clock(clock), .in1(R9466));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9606 (.out1(R9607), .clock(clock), .in1(R9606));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9741 (.out1(R9742), .clock(clock), .in1(R9741));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9923 (.out1(R9924), .clock(clock), .in1(R9923));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10050 (.out1(R10051), .clock(clock), .in1(R10050));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10172 (.out1(R10173), .clock(clock), .in1(R10172));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10341 (.out1(R10342), .clock(clock), .in1(R10341));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10454 (.out1(R10455), .clock(clock), .in1(R10454));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10562 (.out1(R10563), .clock(clock), .in1(R10562));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10718 (.out1(R10719), .clock(clock), .in1(R10718));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10818 (.out1(R10819), .clock(clock), .in1(R10818));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10913 (.out1(R10914), .clock(clock), .in1(R10913));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11055 (.out1(R11056), .clock(clock), .in1(R11055));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11142 (.out1(R11143), .clock(clock), .in1(R11142));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11224 (.out1(R11225), .clock(clock), .in1(R11224));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11353 (.out1(R11354), .clock(clock), .in1(R11353));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11427 (.out1(R11428), .clock(clock), .in1(R11427));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11496 (.out1(R11497), .clock(clock), .in1(R11496));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11612 (.out1(R11613), .clock(clock), .in1(R11612));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11673 (.out1(R11674), .clock(clock), .in1(R11673));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11729 (.out1(R11730), .clock(clock), .in1(R11729));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11832 (.out1(R11833), .clock(clock), .in1(R11832));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11880 (.out1(R11881), .clock(clock), .in1(_1440));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(5), .BITSIZE_out1(64), .PRECISION(64)) op1482 (.out1(_1435), .in1(ip2_3602_D), .in2(5 'd 16));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1483 (.out1(_1436), .in1(_1435));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op1484 (.out1(off_3659), .in1(_1436), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1489 (.out1(_1441), .in1(R11881), .in2(off_3659));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3889 (.out1(R3890), .clock(clock), .in1(R3889));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4145 (.out1(R4146), .clock(clock), .in1(R4145));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4400 (.out1(R4401), .clock(clock), .in1(R4400));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4645 (.out1(R4646), .clock(clock), .in1(R4645));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4885 (.out1(R4886), .clock(clock), .in1(R4885));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5172 (.out1(R5173), .clock(clock), .in1(R5172));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5404 (.out1(R5405), .clock(clock), .in1(R5404));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5631 (.out1(R5632), .clock(clock), .in1(R5631));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5905 (.out1(R5906), .clock(clock), .in1(R5905));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6123 (.out1(R6124), .clock(clock), .in1(R6123));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6336 (.out1(R6337), .clock(clock), .in1(R6336));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6597 (.out1(R6598), .clock(clock), .in1(R6597));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6802 (.out1(R6803), .clock(clock), .in1(R6802));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7002 (.out1(R7003), .clock(clock), .in1(R7002));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7249 (.out1(R7250), .clock(clock), .in1(R7249));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7441 (.out1(R7442), .clock(clock), .in1(R7441));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7628 (.out1(R7629), .clock(clock), .in1(R7628));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7862 (.out1(R7863), .clock(clock), .in1(R7862));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8041 (.out1(R8042), .clock(clock), .in1(R8041));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8215 (.out1(R8216), .clock(clock), .in1(R8215));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8436 (.out1(R8437), .clock(clock), .in1(R8436));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8602 (.out1(R8603), .clock(clock), .in1(R8602));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8763 (.out1(R8764), .clock(clock), .in1(R8763));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8971 (.out1(R8972), .clock(clock), .in1(R8971));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9124 (.out1(R9125), .clock(clock), .in1(R9124));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9272 (.out1(R9273), .clock(clock), .in1(R9272));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9467 (.out1(R9468), .clock(clock), .in1(R9467));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9607 (.out1(R9608), .clock(clock), .in1(R9607));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9742 (.out1(R9743), .clock(clock), .in1(R9742));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9924 (.out1(R9925), .clock(clock), .in1(R9924));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10051 (.out1(R10052), .clock(clock), .in1(R10051));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10173 (.out1(R10174), .clock(clock), .in1(R10173));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10342 (.out1(R10343), .clock(clock), .in1(R10342));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10455 (.out1(R10456), .clock(clock), .in1(R10455));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10563 (.out1(R10564), .clock(clock), .in1(R10563));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10719 (.out1(R10720), .clock(clock), .in1(R10719));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10819 (.out1(R10820), .clock(clock), .in1(R10819));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10914 (.out1(R10915), .clock(clock), .in1(R10914));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11056 (.out1(R11057), .clock(clock), .in1(R11056));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11143 (.out1(R11144), .clock(clock), .in1(R11143));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11225 (.out1(R11226), .clock(clock), .in1(R11225));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11354 (.out1(R11355), .clock(clock), .in1(R11354));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11428 (.out1(R11429), .clock(clock), .in1(R11428));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11497 (.out1(R11498), .clock(clock), .in1(R11497));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11613 (.out1(R11614), .clock(clock), .in1(R11613));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11674 (.out1(R11675), .clock(clock), .in1(R11674));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11730 (.out1(R11731), .clock(clock), .in1(R11730));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11833 (.out1(R11834), .clock(clock), .in1(R11833));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11881 (.out1(R11882), .clock(clock), .in1(off_3659));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11924 (.out1(R11925), .clock(clock), .in1(_1441));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op1490 (.out1(_1442), .in1(R11925), .in2(1 'd 1));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op1491 (.out1(ifout1491), .in1(_1442), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1559 (.out1(_1510), .in1(R11834));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1552 (.out1(_1503), .in1(R11834));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1541 (.out1(_1492), .in1(R11834));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1521 (.out1(_1472), .in1(R11834));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1560 (.out1(_1511), .in1(_1510), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1553 (.out1(_1504), .in1(_1503), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1542 (.out1(_1493), .in1(_1492), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1522 (.out1(_1473), .in1(_1472), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3890 (.out1(R3891), .clock(clock), .in1(R3890));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4146 (.out1(R4147), .clock(clock), .in1(R4146));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4401 (.out1(R4402), .clock(clock), .in1(R4401));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4646 (.out1(R4647), .clock(clock), .in1(R4646));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4886 (.out1(R4887), .clock(clock), .in1(R4886));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5173 (.out1(R5174), .clock(clock), .in1(R5173));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5405 (.out1(R5406), .clock(clock), .in1(R5405));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5632 (.out1(R5633), .clock(clock), .in1(R5632));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5906 (.out1(R5907), .clock(clock), .in1(R5906));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6124 (.out1(R6125), .clock(clock), .in1(R6124));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6337 (.out1(R6338), .clock(clock), .in1(R6337));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6598 (.out1(R6599), .clock(clock), .in1(R6598));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6803 (.out1(R6804), .clock(clock), .in1(R6803));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7003 (.out1(R7004), .clock(clock), .in1(R7003));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7250 (.out1(R7251), .clock(clock), .in1(R7250));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7442 (.out1(R7443), .clock(clock), .in1(R7442));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7629 (.out1(R7630), .clock(clock), .in1(R7629));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7863 (.out1(R7864), .clock(clock), .in1(R7863));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8042 (.out1(R8043), .clock(clock), .in1(R8042));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8216 (.out1(R8217), .clock(clock), .in1(R8216));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8437 (.out1(R8438), .clock(clock), .in1(R8437));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8603 (.out1(R8604), .clock(clock), .in1(R8603));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8764 (.out1(R8765), .clock(clock), .in1(R8764));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8972 (.out1(R8973), .clock(clock), .in1(R8972));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9125 (.out1(R9126), .clock(clock), .in1(R9125));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9273 (.out1(R9274), .clock(clock), .in1(R9273));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9468 (.out1(R9469), .clock(clock), .in1(R9468));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9608 (.out1(R9609), .clock(clock), .in1(R9608));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9743 (.out1(R9744), .clock(clock), .in1(R9743));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9925 (.out1(R9926), .clock(clock), .in1(R9925));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10052 (.out1(R10053), .clock(clock), .in1(R10052));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10174 (.out1(R10175), .clock(clock), .in1(R10174));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10343 (.out1(R10344), .clock(clock), .in1(R10343));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10456 (.out1(R10457), .clock(clock), .in1(R10456));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10564 (.out1(R10565), .clock(clock), .in1(R10564));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10720 (.out1(R10721), .clock(clock), .in1(R10720));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10820 (.out1(R10821), .clock(clock), .in1(R10820));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10915 (.out1(R10916), .clock(clock), .in1(R10915));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11057 (.out1(R11058), .clock(clock), .in1(R11057));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11144 (.out1(R11145), .clock(clock), .in1(R11144));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11226 (.out1(R11227), .clock(clock), .in1(R11226));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11355 (.out1(R11356), .clock(clock), .in1(R11355));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11429 (.out1(R11430), .clock(clock), .in1(R11429));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11498 (.out1(R11499), .clock(clock), .in1(R11498));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11614 (.out1(R11615), .clock(clock), .in1(R11614));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11675 (.out1(R11676), .clock(clock), .in1(R11675));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11731 (.out1(R11732), .clock(clock), .in1(R11731));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11834 (.out1(R11835), .clock(clock), .in1(R11834));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11882 (.out1(R11883), .clock(clock), .in1(R11882));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11925 (.out1(R11926), .clock(clock), .in1(ifout1491));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11975 (.out1(R11976), .clock(clock), .in1(_1511));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11976 (.out1(R11977), .clock(clock), .in1(_1504));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11977 (.out1(R11978), .clock(clock), .in1(_1493));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11978 (.out1(R11979), .clock(clock), .in1(_1473));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1534 (.out1(_1485), .in1(R11835));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1514 (.out1(_1465), .in1(R11835));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1503 (.out1(_1454), .in1(R11835));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1496 (.out1(_1447), .in1(R11835));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1563 (.out1(_1514), .in1(2 'd 2), .in2(R11883));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1535 (.out1(_1486), .in1(_1485), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1515 (.out1(_1466), .in1(_1465), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1504 (.out1(_1455), .in1(_1454), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1497 (.out1(_1448), .in1(_1447), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1561 (.out1(_1512), .in1(vec106_3660_D), .in2(R11976));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1554 (.out1(_1505), .in1(vec106_3660_D), .in2(R11977));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1543 (.out1(_1494), .in1(vec106_3660_D), .in2(R11978));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1523 (.out1(_1474), .in1(vec106_3660_D), .in2(R11979));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3891 (.out1(R3892), .clock(clock), .in1(R3891));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4147 (.out1(R4148), .clock(clock), .in1(R4147));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4402 (.out1(R4403), .clock(clock), .in1(R4402));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4647 (.out1(R4648), .clock(clock), .in1(R4647));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4887 (.out1(R4888), .clock(clock), .in1(R4887));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5174 (.out1(R5175), .clock(clock), .in1(R5174));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5406 (.out1(R5407), .clock(clock), .in1(R5406));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5633 (.out1(R5634), .clock(clock), .in1(R5633));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5907 (.out1(R5908), .clock(clock), .in1(R5907));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6125 (.out1(R6126), .clock(clock), .in1(R6125));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6338 (.out1(R6339), .clock(clock), .in1(R6338));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6599 (.out1(R6600), .clock(clock), .in1(R6599));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6804 (.out1(R6805), .clock(clock), .in1(R6804));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7004 (.out1(R7005), .clock(clock), .in1(R7004));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7251 (.out1(R7252), .clock(clock), .in1(R7251));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7443 (.out1(R7444), .clock(clock), .in1(R7443));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7630 (.out1(R7631), .clock(clock), .in1(R7630));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7864 (.out1(R7865), .clock(clock), .in1(R7864));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8043 (.out1(R8044), .clock(clock), .in1(R8043));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8217 (.out1(R8218), .clock(clock), .in1(R8217));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8438 (.out1(R8439), .clock(clock), .in1(R8438));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8604 (.out1(R8605), .clock(clock), .in1(R8604));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8765 (.out1(R8766), .clock(clock), .in1(R8765));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8973 (.out1(R8974), .clock(clock), .in1(R8973));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9126 (.out1(R9127), .clock(clock), .in1(R9126));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9274 (.out1(R9275), .clock(clock), .in1(R9274));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9469 (.out1(R9470), .clock(clock), .in1(R9469));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9609 (.out1(R9610), .clock(clock), .in1(R9609));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9744 (.out1(R9745), .clock(clock), .in1(R9744));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9926 (.out1(R9927), .clock(clock), .in1(R9926));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10053 (.out1(R10054), .clock(clock), .in1(R10053));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10175 (.out1(R10176), .clock(clock), .in1(R10175));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10344 (.out1(R10345), .clock(clock), .in1(R10344));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10457 (.out1(R10458), .clock(clock), .in1(R10457));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10565 (.out1(R10566), .clock(clock), .in1(R10565));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10721 (.out1(R10722), .clock(clock), .in1(R10721));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10821 (.out1(R10822), .clock(clock), .in1(R10821));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10916 (.out1(R10917), .clock(clock), .in1(R10916));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11058 (.out1(R11059), .clock(clock), .in1(R11058));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11145 (.out1(R11146), .clock(clock), .in1(R11145));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11227 (.out1(R11228), .clock(clock), .in1(R11227));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11356 (.out1(R11357), .clock(clock), .in1(R11356));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11430 (.out1(R11431), .clock(clock), .in1(R11430));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11499 (.out1(R11500), .clock(clock), .in1(R11499));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11615 (.out1(R11616), .clock(clock), .in1(R11615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11676 (.out1(R11677), .clock(clock), .in1(R11676));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11732 (.out1(R11733), .clock(clock), .in1(R11732));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11835 (.out1(R11836), .clock(clock), .in1(R11835));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11883 (.out1(R11884), .clock(clock), .in1(R11883));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11926 (.out1(R11927), .clock(clock), .in1(R11926));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11979 (.out1(R11980), .clock(clock), .in1(_1514));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11980 (.out1(R11981), .clock(clock), .in1(_1486));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11981 (.out1(R11982), .clock(clock), .in1(_1466));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11982 (.out1(R11983), .clock(clock), .in1(_1455));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11983 (.out1(R11984), .clock(clock), .in1(_1448));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11984 (.out1(R11985), .clock(clock), .in1(_1512));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11985 (.out1(R11986), .clock(clock), .in1(_1505));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11986 (.out1(R11987), .clock(clock), .in1(_1494));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11987 (.out1(R11988), .clock(clock), .in1(_1474));
  SRAM op1562 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1513),.ADR(R11985));
  SRAM op1555 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1506),.ADR(R11986));
  SRAM op1544 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1495),.ADR(R11987));
  SRAM op1524 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1475),.ADR(R11988));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1556 (.out1(_1507), .in1(2 'd 2), .in2(R11884));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1545 (.out1(_1496), .in1(2 'd 2), .in2(R11884));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1538 (.out1(_1489), .in1(2 'd 2), .in2(R11884));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1525 (.out1(_1476), .in1(2 'd 2), .in2(R11884));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1518 (.out1(_1469), .in1(2 'd 2), .in2(R11884));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1507 (.out1(_1458), .in1(2 'd 2), .in2(R11884));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1536 (.out1(_1487), .in1(vec106_3660_D), .in2(R11981));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1516 (.out1(_1467), .in1(vec106_3660_D), .in2(R11982));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1505 (.out1(_1456), .in1(vec106_3660_D), .in2(R11983));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1498 (.out1(_1449), .in1(vec106_3660_D), .in2(R11984));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1564 (.out1(_1515), .in1(R11980), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3892 (.out1(R3893), .clock(clock), .in1(R3892));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4148 (.out1(R4149), .clock(clock), .in1(R4148));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4403 (.out1(R4404), .clock(clock), .in1(R4403));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4648 (.out1(R4649), .clock(clock), .in1(R4648));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4888 (.out1(R4889), .clock(clock), .in1(R4888));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5175 (.out1(R5176), .clock(clock), .in1(R5175));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5407 (.out1(R5408), .clock(clock), .in1(R5407));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5634 (.out1(R5635), .clock(clock), .in1(R5634));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5908 (.out1(R5909), .clock(clock), .in1(R5908));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6126 (.out1(R6127), .clock(clock), .in1(R6126));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6339 (.out1(R6340), .clock(clock), .in1(R6339));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6600 (.out1(R6601), .clock(clock), .in1(R6600));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6805 (.out1(R6806), .clock(clock), .in1(R6805));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7005 (.out1(R7006), .clock(clock), .in1(R7005));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7252 (.out1(R7253), .clock(clock), .in1(R7252));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7444 (.out1(R7445), .clock(clock), .in1(R7444));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7631 (.out1(R7632), .clock(clock), .in1(R7631));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7865 (.out1(R7866), .clock(clock), .in1(R7865));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8044 (.out1(R8045), .clock(clock), .in1(R8044));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8218 (.out1(R8219), .clock(clock), .in1(R8218));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8439 (.out1(R8440), .clock(clock), .in1(R8439));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8605 (.out1(R8606), .clock(clock), .in1(R8605));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8766 (.out1(R8767), .clock(clock), .in1(R8766));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8974 (.out1(R8975), .clock(clock), .in1(R8974));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9127 (.out1(R9128), .clock(clock), .in1(R9127));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9275 (.out1(R9276), .clock(clock), .in1(R9275));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9470 (.out1(R9471), .clock(clock), .in1(R9470));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9610 (.out1(R9611), .clock(clock), .in1(R9610));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9745 (.out1(R9746), .clock(clock), .in1(R9745));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9927 (.out1(R9928), .clock(clock), .in1(R9927));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10054 (.out1(R10055), .clock(clock), .in1(R10054));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10176 (.out1(R10177), .clock(clock), .in1(R10176));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10345 (.out1(R10346), .clock(clock), .in1(R10345));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10458 (.out1(R10459), .clock(clock), .in1(R10458));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10566 (.out1(R10567), .clock(clock), .in1(R10566));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10722 (.out1(R10723), .clock(clock), .in1(R10722));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10822 (.out1(R10823), .clock(clock), .in1(R10822));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10917 (.out1(R10918), .clock(clock), .in1(R10917));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11059 (.out1(R11060), .clock(clock), .in1(R11059));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11146 (.out1(R11147), .clock(clock), .in1(R11146));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11228 (.out1(R11229), .clock(clock), .in1(R11228));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11357 (.out1(R11358), .clock(clock), .in1(R11357));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11431 (.out1(R11432), .clock(clock), .in1(R11431));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11500 (.out1(R11501), .clock(clock), .in1(R11500));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11616 (.out1(R11617), .clock(clock), .in1(R11616));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11677 (.out1(R11678), .clock(clock), .in1(R11677));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11733 (.out1(R11734), .clock(clock), .in1(R11733));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11836 (.out1(R11837), .clock(clock), .in1(R11836));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11884 (.out1(R11885), .clock(clock), .in1(R11884));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11927 (.out1(R11928), .clock(clock), .in1(R11927));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11988 (.out1(R11989), .clock(clock), .in1(_1513));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11989 (.out1(R11990), .clock(clock), .in1(_1506));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11990 (.out1(R11991), .clock(clock), .in1(_1495));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11991 (.out1(R11992), .clock(clock), .in1(_1475));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11992 (.out1(R11993), .clock(clock), .in1(_1507));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11993 (.out1(R11994), .clock(clock), .in1(_1496));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11994 (.out1(R11995), .clock(clock), .in1(_1489));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11995 (.out1(R11996), .clock(clock), .in1(_1476));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11996 (.out1(R11997), .clock(clock), .in1(_1469));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11997 (.out1(R11998), .clock(clock), .in1(_1458));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11998 (.out1(R11999), .clock(clock), .in1(_1487));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op11999 (.out1(R12000), .clock(clock), .in1(_1467));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12000 (.out1(R12001), .clock(clock), .in1(_1456));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12001 (.out1(R12002), .clock(clock), .in1(_1449));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12002 (.out1(R12003), .clock(clock), .in1(_1515));
  SRAM op1537 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1488),.ADR(R11999));
  SRAM op1517 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1468),.ADR(R12000));
  SRAM op1506 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1457),.ADR(R12001));
  SRAM op1499 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1450),.ADR(R12002));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1565 (.out1(_1516), .in1(R11989), .in2(R12003));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1566 (.out1(_1517), .in1(_1516), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1557 (.out1(_1508), .in1(R11993), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1546 (.out1(_1497), .in1(R11994), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1526 (.out1(_1477), .in1(R11996), .in2(64 'd 18446744073709551615));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1500 (.out1(_1451), .in1(2 'd 2), .in2(R11885));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1567 (.out1(_1518), .in1(_1517), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1558 (.out1(_1509), .in1(R11990), .in2(_1508));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1547 (.out1(_1498), .in1(R11991), .in2(_1497));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1527 (.out1(_1478), .in1(R11992), .in2(_1477));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1568 (.out1(_1519), .in1(_1509), .in2(_1518));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1548 (.out1(_1499), .in1(_1498), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1539 (.out1(_1490), .in1(R11995), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1528 (.out1(_1479), .in1(_1478), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1519 (.out1(_1470), .in1(R11997), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1508 (.out1(_1459), .in1(R11998), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3893 (.out1(R3894), .clock(clock), .in1(R3893));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4149 (.out1(R4150), .clock(clock), .in1(R4149));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4404 (.out1(R4405), .clock(clock), .in1(R4404));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4649 (.out1(R4650), .clock(clock), .in1(R4649));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4889 (.out1(R4890), .clock(clock), .in1(R4889));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5176 (.out1(R5177), .clock(clock), .in1(R5176));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5408 (.out1(R5409), .clock(clock), .in1(R5408));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5635 (.out1(R5636), .clock(clock), .in1(R5635));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5909 (.out1(R5910), .clock(clock), .in1(R5909));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6127 (.out1(R6128), .clock(clock), .in1(R6127));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6340 (.out1(R6341), .clock(clock), .in1(R6340));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6601 (.out1(R6602), .clock(clock), .in1(R6601));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6806 (.out1(R6807), .clock(clock), .in1(R6806));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7006 (.out1(R7007), .clock(clock), .in1(R7006));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7253 (.out1(R7254), .clock(clock), .in1(R7253));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7445 (.out1(R7446), .clock(clock), .in1(R7445));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7632 (.out1(R7633), .clock(clock), .in1(R7632));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7866 (.out1(R7867), .clock(clock), .in1(R7866));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8045 (.out1(R8046), .clock(clock), .in1(R8045));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8219 (.out1(R8220), .clock(clock), .in1(R8219));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8440 (.out1(R8441), .clock(clock), .in1(R8440));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8606 (.out1(R8607), .clock(clock), .in1(R8606));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8767 (.out1(R8768), .clock(clock), .in1(R8767));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8975 (.out1(R8976), .clock(clock), .in1(R8975));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9128 (.out1(R9129), .clock(clock), .in1(R9128));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9276 (.out1(R9277), .clock(clock), .in1(R9276));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9471 (.out1(R9472), .clock(clock), .in1(R9471));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9611 (.out1(R9612), .clock(clock), .in1(R9611));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9746 (.out1(R9747), .clock(clock), .in1(R9746));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9928 (.out1(R9929), .clock(clock), .in1(R9928));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10055 (.out1(R10056), .clock(clock), .in1(R10055));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10177 (.out1(R10178), .clock(clock), .in1(R10177));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10346 (.out1(R10347), .clock(clock), .in1(R10346));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10459 (.out1(R10460), .clock(clock), .in1(R10459));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10567 (.out1(R10568), .clock(clock), .in1(R10567));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10723 (.out1(R10724), .clock(clock), .in1(R10723));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10823 (.out1(R10824), .clock(clock), .in1(R10823));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10918 (.out1(R10919), .clock(clock), .in1(R10918));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11060 (.out1(R11061), .clock(clock), .in1(R11060));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11147 (.out1(R11148), .clock(clock), .in1(R11147));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11229 (.out1(R11230), .clock(clock), .in1(R11229));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11358 (.out1(R11359), .clock(clock), .in1(R11358));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11432 (.out1(R11433), .clock(clock), .in1(R11432));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11501 (.out1(R11502), .clock(clock), .in1(R11501));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11617 (.out1(R11618), .clock(clock), .in1(R11617));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11678 (.out1(R11679), .clock(clock), .in1(R11678));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11734 (.out1(R11735), .clock(clock), .in1(R11734));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11837 (.out1(R11838), .clock(clock), .in1(R11837));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11885 (.out1(R11886), .clock(clock), .in1(R11885));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11928 (.out1(R11929), .clock(clock), .in1(R11928));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12003 (.out1(R12004), .clock(clock), .in1(_1488));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12004 (.out1(R12005), .clock(clock), .in1(_1468));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12005 (.out1(R12006), .clock(clock), .in1(_1457));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12006 (.out1(R12007), .clock(clock), .in1(_1450));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12007 (.out1(R12008), .clock(clock), .in1(_1451));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12008 (.out1(R12009), .clock(clock), .in1(_1519));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12009 (.out1(R12010), .clock(clock), .in1(_1499));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12010 (.out1(R12011), .clock(clock), .in1(_1490));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12011 (.out1(R12012), .clock(clock), .in1(_1479));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12012 (.out1(R12013), .clock(clock), .in1(_1470));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12013 (.out1(R12014), .clock(clock), .in1(_1459));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1549 (.out1(_1500), .in1(R12010), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1540 (.out1(_1491), .in1(R12004), .in2(R12011));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1509 (.out1(_1460), .in1(R12006), .in2(R12014));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1569 (.out1(_1520), .in1(R12009), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1550 (.out1(_1501), .in1(_1491), .in2(_1500));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1529 (.out1(_1480), .in1(R12012), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1520 (.out1(_1471), .in1(R12005), .in2(R12013));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1510 (.out1(_1461), .in1(_1460), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1501 (.out1(_1452), .in1(R12008), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1530 (.out1(_1481), .in1(_1471), .in2(_1480));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1570 (.out1(_1521), .in1(_1520), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1551 (.out1(_1502), .in1(_1501), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1511 (.out1(_1462), .in1(_1461), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1502 (.out1(_1453), .in1(R12007), .in2(_1452));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1571 (.out1(_1522), .in1(_1502), .in2(_1521));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1531 (.out1(_1482), .in1(_1481), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1512 (.out1(_1463), .in1(_1453), .in2(_1462));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3894 (.out1(R3895), .clock(clock), .in1(R3894));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4150 (.out1(R4151), .clock(clock), .in1(R4150));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4405 (.out1(R4406), .clock(clock), .in1(R4405));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4650 (.out1(R4651), .clock(clock), .in1(R4650));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4890 (.out1(R4891), .clock(clock), .in1(R4890));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5177 (.out1(R5178), .clock(clock), .in1(R5177));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5409 (.out1(R5410), .clock(clock), .in1(R5409));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5636 (.out1(R5637), .clock(clock), .in1(R5636));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5910 (.out1(R5911), .clock(clock), .in1(R5910));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6128 (.out1(R6129), .clock(clock), .in1(R6128));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6341 (.out1(R6342), .clock(clock), .in1(R6341));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6602 (.out1(R6603), .clock(clock), .in1(R6602));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6807 (.out1(R6808), .clock(clock), .in1(R6807));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7007 (.out1(R7008), .clock(clock), .in1(R7007));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7254 (.out1(R7255), .clock(clock), .in1(R7254));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7446 (.out1(R7447), .clock(clock), .in1(R7446));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7633 (.out1(R7634), .clock(clock), .in1(R7633));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7867 (.out1(R7868), .clock(clock), .in1(R7867));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8046 (.out1(R8047), .clock(clock), .in1(R8046));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8220 (.out1(R8221), .clock(clock), .in1(R8220));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8441 (.out1(R8442), .clock(clock), .in1(R8441));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8607 (.out1(R8608), .clock(clock), .in1(R8607));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8768 (.out1(R8769), .clock(clock), .in1(R8768));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8976 (.out1(R8977), .clock(clock), .in1(R8976));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9129 (.out1(R9130), .clock(clock), .in1(R9129));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9277 (.out1(R9278), .clock(clock), .in1(R9277));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9472 (.out1(R9473), .clock(clock), .in1(R9472));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9612 (.out1(R9613), .clock(clock), .in1(R9612));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9747 (.out1(R9748), .clock(clock), .in1(R9747));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9929 (.out1(R9930), .clock(clock), .in1(R9929));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10056 (.out1(R10057), .clock(clock), .in1(R10056));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10178 (.out1(R10179), .clock(clock), .in1(R10178));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10347 (.out1(R10348), .clock(clock), .in1(R10347));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10460 (.out1(R10461), .clock(clock), .in1(R10460));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10568 (.out1(R10569), .clock(clock), .in1(R10568));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10724 (.out1(R10725), .clock(clock), .in1(R10724));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10824 (.out1(R10825), .clock(clock), .in1(R10824));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10919 (.out1(R10920), .clock(clock), .in1(R10919));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11061 (.out1(R11062), .clock(clock), .in1(R11061));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11148 (.out1(R11149), .clock(clock), .in1(R11148));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11230 (.out1(R11231), .clock(clock), .in1(R11230));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11359 (.out1(R11360), .clock(clock), .in1(R11359));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11433 (.out1(R11434), .clock(clock), .in1(R11433));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11502 (.out1(R11503), .clock(clock), .in1(R11502));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11618 (.out1(R11619), .clock(clock), .in1(R11618));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11679 (.out1(R11680), .clock(clock), .in1(R11679));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11735 (.out1(R11736), .clock(clock), .in1(R11735));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11838 (.out1(R11839), .clock(clock), .in1(R11838));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11886 (.out1(R11887), .clock(clock), .in1(R11886));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11929 (.out1(R11930), .clock(clock), .in1(R11929));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12014 (.out1(R12015), .clock(clock), .in1(_1522));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12015 (.out1(R12016), .clock(clock), .in1(_1482));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12016 (.out1(R12017), .clock(clock), .in1(_1463));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1492 (.out1(_1443), .in1(R11839));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1532 (.out1(_1483), .in1(R12016), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1513 (.out1(_1464), .in1(R12017), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op1572 (.out1(_1523), .in1(R12015), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1533 (.out1(_1484), .in1(_1464), .in2(_1483));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1493 (.out1(_1444), .in1(_1443), .in2(2 'd 2));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1573 (.out1(_1524), .in1(_1484), .in2(_1523));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op1574 (.out1(_1525), .in1(_1524), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3895 (.out1(R3896), .clock(clock), .in1(R3895));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4151 (.out1(R4152), .clock(clock), .in1(R4151));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4406 (.out1(R4407), .clock(clock), .in1(R4406));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4651 (.out1(R4652), .clock(clock), .in1(R4651));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4891 (.out1(R4892), .clock(clock), .in1(R4891));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5178 (.out1(R5179), .clock(clock), .in1(R5178));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5410 (.out1(R5411), .clock(clock), .in1(R5410));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5637 (.out1(R5638), .clock(clock), .in1(R5637));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5911 (.out1(R5912), .clock(clock), .in1(R5911));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6129 (.out1(R6130), .clock(clock), .in1(R6129));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6342 (.out1(R6343), .clock(clock), .in1(R6342));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6603 (.out1(R6604), .clock(clock), .in1(R6603));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6808 (.out1(R6809), .clock(clock), .in1(R6808));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7008 (.out1(R7009), .clock(clock), .in1(R7008));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7255 (.out1(R7256), .clock(clock), .in1(R7255));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7447 (.out1(R7448), .clock(clock), .in1(R7447));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7634 (.out1(R7635), .clock(clock), .in1(R7634));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7868 (.out1(R7869), .clock(clock), .in1(R7868));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8047 (.out1(R8048), .clock(clock), .in1(R8047));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8221 (.out1(R8222), .clock(clock), .in1(R8221));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8442 (.out1(R8443), .clock(clock), .in1(R8442));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8608 (.out1(R8609), .clock(clock), .in1(R8608));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8769 (.out1(R8770), .clock(clock), .in1(R8769));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8977 (.out1(R8978), .clock(clock), .in1(R8977));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9130 (.out1(R9131), .clock(clock), .in1(R9130));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9278 (.out1(R9279), .clock(clock), .in1(R9278));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9473 (.out1(R9474), .clock(clock), .in1(R9473));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9613 (.out1(R9614), .clock(clock), .in1(R9613));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9748 (.out1(R9749), .clock(clock), .in1(R9748));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9930 (.out1(R9931), .clock(clock), .in1(R9930));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10057 (.out1(R10058), .clock(clock), .in1(R10057));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10179 (.out1(R10180), .clock(clock), .in1(R10179));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10348 (.out1(R10349), .clock(clock), .in1(R10348));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10461 (.out1(R10462), .clock(clock), .in1(R10461));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10569 (.out1(R10570), .clock(clock), .in1(R10569));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10725 (.out1(R10726), .clock(clock), .in1(R10725));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10825 (.out1(R10826), .clock(clock), .in1(R10825));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10920 (.out1(R10921), .clock(clock), .in1(R10920));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11062 (.out1(R11063), .clock(clock), .in1(R11062));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11149 (.out1(R11150), .clock(clock), .in1(R11149));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11231 (.out1(R11232), .clock(clock), .in1(R11231));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11360 (.out1(R11361), .clock(clock), .in1(R11360));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11434 (.out1(R11435), .clock(clock), .in1(R11434));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11503 (.out1(R11504), .clock(clock), .in1(R11503));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11619 (.out1(R11620), .clock(clock), .in1(R11619));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11680 (.out1(R11681), .clock(clock), .in1(R11680));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11736 (.out1(R11737), .clock(clock), .in1(R11736));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11839 (.out1(R11840), .clock(clock), .in1(R11839));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11887 (.out1(R11888), .clock(clock), .in1(R11887));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11930 (.out1(R11931), .clock(clock), .in1(R11930));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12017 (.out1(R12018), .clock(clock), .in1(_1444));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12018 (.out1(R12019), .clock(clock), .in1(_1525));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op1575 (.out1(_1526), .in1(R12019), .in2(57 'd 72340172838076673));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1494 (.out1(_1445), .in1(base0_106_3665_D), .in2(R12018));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3896 (.out1(R3897), .clock(clock), .in1(R3896));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4152 (.out1(R4153), .clock(clock), .in1(R4152));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4407 (.out1(R4408), .clock(clock), .in1(R4407));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4652 (.out1(R4653), .clock(clock), .in1(R4652));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4892 (.out1(R4893), .clock(clock), .in1(R4892));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5179 (.out1(R5180), .clock(clock), .in1(R5179));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5411 (.out1(R5412), .clock(clock), .in1(R5411));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5638 (.out1(R5639), .clock(clock), .in1(R5638));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5912 (.out1(R5913), .clock(clock), .in1(R5912));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6130 (.out1(R6131), .clock(clock), .in1(R6130));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6343 (.out1(R6344), .clock(clock), .in1(R6343));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6604 (.out1(R6605), .clock(clock), .in1(R6604));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6809 (.out1(R6810), .clock(clock), .in1(R6809));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7009 (.out1(R7010), .clock(clock), .in1(R7009));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7256 (.out1(R7257), .clock(clock), .in1(R7256));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7448 (.out1(R7449), .clock(clock), .in1(R7448));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7635 (.out1(R7636), .clock(clock), .in1(R7635));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7869 (.out1(R7870), .clock(clock), .in1(R7869));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8048 (.out1(R8049), .clock(clock), .in1(R8048));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8222 (.out1(R8223), .clock(clock), .in1(R8222));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8443 (.out1(R8444), .clock(clock), .in1(R8443));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8609 (.out1(R8610), .clock(clock), .in1(R8609));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8770 (.out1(R8771), .clock(clock), .in1(R8770));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8978 (.out1(R8979), .clock(clock), .in1(R8978));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9131 (.out1(R9132), .clock(clock), .in1(R9131));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9279 (.out1(R9280), .clock(clock), .in1(R9279));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9474 (.out1(R9475), .clock(clock), .in1(R9474));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9614 (.out1(R9615), .clock(clock), .in1(R9614));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9749 (.out1(R9750), .clock(clock), .in1(R9749));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9931 (.out1(R9932), .clock(clock), .in1(R9931));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10058 (.out1(R10059), .clock(clock), .in1(R10058));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10180 (.out1(R10181), .clock(clock), .in1(R10180));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10349 (.out1(R10350), .clock(clock), .in1(R10349));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10462 (.out1(R10463), .clock(clock), .in1(R10462));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10570 (.out1(R10571), .clock(clock), .in1(R10570));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10726 (.out1(R10727), .clock(clock), .in1(R10726));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10826 (.out1(R10827), .clock(clock), .in1(R10826));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10921 (.out1(R10922), .clock(clock), .in1(R10921));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11063 (.out1(R11064), .clock(clock), .in1(R11063));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11150 (.out1(R11151), .clock(clock), .in1(R11150));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11232 (.out1(R11233), .clock(clock), .in1(R11232));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11361 (.out1(R11362), .clock(clock), .in1(R11361));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11435 (.out1(R11436), .clock(clock), .in1(R11435));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11504 (.out1(R11505), .clock(clock), .in1(R11504));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11620 (.out1(R11621), .clock(clock), .in1(R11620));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11681 (.out1(R11682), .clock(clock), .in1(R11681));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11737 (.out1(R11738), .clock(clock), .in1(R11737));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11840 (.out1(R11841), .clock(clock), .in1(R11840));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11888 (.out1(R11889), .clock(clock), .in1(R11888));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11931 (.out1(R11932), .clock(clock), .in1(R11931));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12019 (.out1(R12020), .clock(clock), .in1(_1526));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12020 (.out1(R12021), .clock(clock), .in1(_1445));
  SRAM op1495 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1446),.ADR(R12021));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op1576 (.out1(_1527), .in1(R12020), .in2(6 'd 56));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3897 (.out1(R3898), .clock(clock), .in1(R3897));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4153 (.out1(R4154), .clock(clock), .in1(R4153));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4408 (.out1(R4409), .clock(clock), .in1(R4408));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4653 (.out1(R4654), .clock(clock), .in1(R4653));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4893 (.out1(R4894), .clock(clock), .in1(R4893));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5180 (.out1(R5181), .clock(clock), .in1(R5180));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5412 (.out1(R5413), .clock(clock), .in1(R5412));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5639 (.out1(R5640), .clock(clock), .in1(R5639));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5913 (.out1(R5914), .clock(clock), .in1(R5913));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6131 (.out1(R6132), .clock(clock), .in1(R6131));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6344 (.out1(R6345), .clock(clock), .in1(R6344));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6605 (.out1(R6606), .clock(clock), .in1(R6605));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6810 (.out1(R6811), .clock(clock), .in1(R6810));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7010 (.out1(R7011), .clock(clock), .in1(R7010));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7257 (.out1(R7258), .clock(clock), .in1(R7257));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7449 (.out1(R7450), .clock(clock), .in1(R7449));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7636 (.out1(R7637), .clock(clock), .in1(R7636));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7870 (.out1(R7871), .clock(clock), .in1(R7870));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8049 (.out1(R8050), .clock(clock), .in1(R8049));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8223 (.out1(R8224), .clock(clock), .in1(R8223));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8444 (.out1(R8445), .clock(clock), .in1(R8444));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8610 (.out1(R8611), .clock(clock), .in1(R8610));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8771 (.out1(R8772), .clock(clock), .in1(R8771));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8979 (.out1(R8980), .clock(clock), .in1(R8979));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9132 (.out1(R9133), .clock(clock), .in1(R9132));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9280 (.out1(R9281), .clock(clock), .in1(R9280));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9475 (.out1(R9476), .clock(clock), .in1(R9475));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9615 (.out1(R9616), .clock(clock), .in1(R9615));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9750 (.out1(R9751), .clock(clock), .in1(R9750));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9932 (.out1(R9933), .clock(clock), .in1(R9932));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10059 (.out1(R10060), .clock(clock), .in1(R10059));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10181 (.out1(R10182), .clock(clock), .in1(R10181));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10350 (.out1(R10351), .clock(clock), .in1(R10350));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10463 (.out1(R10464), .clock(clock), .in1(R10463));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10571 (.out1(R10572), .clock(clock), .in1(R10571));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10727 (.out1(R10728), .clock(clock), .in1(R10727));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10827 (.out1(R10828), .clock(clock), .in1(R10827));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10922 (.out1(R10923), .clock(clock), .in1(R10922));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11064 (.out1(R11065), .clock(clock), .in1(R11064));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11151 (.out1(R11152), .clock(clock), .in1(R11151));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11233 (.out1(R11234), .clock(clock), .in1(R11233));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11362 (.out1(R11363), .clock(clock), .in1(R11362));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11436 (.out1(R11437), .clock(clock), .in1(R11436));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11505 (.out1(R11506), .clock(clock), .in1(R11505));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11621 (.out1(R11622), .clock(clock), .in1(R11621));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11682 (.out1(R11683), .clock(clock), .in1(R11682));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11738 (.out1(R11739), .clock(clock), .in1(R11738));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11841 (.out1(R11842), .clock(clock), .in1(R11841));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11889 (.out1(R11890), .clock(clock), .in1(R11889));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11932 (.out1(R11933), .clock(clock), .in1(R11932));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12021 (.out1(R12022), .clock(clock), .in1(_1446));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12022 (.out1(R12023), .clock(clock), .in1(_1527));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1577 (.out1(_1528), .in1(R12023));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1578 (.out1(_1529), .in1(R12022), .in2(_1528));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1579 (.out1(idx_3666), .in1(_1529), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3898 (.out1(R3899), .clock(clock), .in1(R3898));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4154 (.out1(R4155), .clock(clock), .in1(R4154));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4409 (.out1(R4410), .clock(clock), .in1(R4409));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4654 (.out1(R4655), .clock(clock), .in1(R4654));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4894 (.out1(R4895), .clock(clock), .in1(R4894));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5181 (.out1(R5182), .clock(clock), .in1(R5181));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5413 (.out1(R5414), .clock(clock), .in1(R5413));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5640 (.out1(R5641), .clock(clock), .in1(R5640));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5914 (.out1(R5915), .clock(clock), .in1(R5914));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6132 (.out1(R6133), .clock(clock), .in1(R6132));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6345 (.out1(R6346), .clock(clock), .in1(R6345));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6606 (.out1(R6607), .clock(clock), .in1(R6606));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6811 (.out1(R6812), .clock(clock), .in1(R6811));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7011 (.out1(R7012), .clock(clock), .in1(R7011));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7258 (.out1(R7259), .clock(clock), .in1(R7258));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7450 (.out1(R7451), .clock(clock), .in1(R7450));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7637 (.out1(R7638), .clock(clock), .in1(R7637));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7871 (.out1(R7872), .clock(clock), .in1(R7871));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8050 (.out1(R8051), .clock(clock), .in1(R8050));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8224 (.out1(R8225), .clock(clock), .in1(R8224));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8445 (.out1(R8446), .clock(clock), .in1(R8445));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8611 (.out1(R8612), .clock(clock), .in1(R8611));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8772 (.out1(R8773), .clock(clock), .in1(R8772));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8980 (.out1(R8981), .clock(clock), .in1(R8980));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9133 (.out1(R9134), .clock(clock), .in1(R9133));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9281 (.out1(R9282), .clock(clock), .in1(R9281));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9476 (.out1(R9477), .clock(clock), .in1(R9476));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9616 (.out1(R9617), .clock(clock), .in1(R9616));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9751 (.out1(R9752), .clock(clock), .in1(R9751));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9933 (.out1(R9934), .clock(clock), .in1(R9933));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10060 (.out1(R10061), .clock(clock), .in1(R10060));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10182 (.out1(R10183), .clock(clock), .in1(R10182));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10351 (.out1(R10352), .clock(clock), .in1(R10351));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10464 (.out1(R10465), .clock(clock), .in1(R10464));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10572 (.out1(R10573), .clock(clock), .in1(R10572));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10728 (.out1(R10729), .clock(clock), .in1(R10728));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10828 (.out1(R10829), .clock(clock), .in1(R10828));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10923 (.out1(R10924), .clock(clock), .in1(R10923));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11065 (.out1(R11066), .clock(clock), .in1(R11065));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11152 (.out1(R11153), .clock(clock), .in1(R11152));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11234 (.out1(R11235), .clock(clock), .in1(R11234));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11363 (.out1(R11364), .clock(clock), .in1(R11363));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11437 (.out1(R11438), .clock(clock), .in1(R11437));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11506 (.out1(R11507), .clock(clock), .in1(R11506));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11622 (.out1(R11623), .clock(clock), .in1(R11622));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11683 (.out1(R11684), .clock(clock), .in1(R11683));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11739 (.out1(R11740), .clock(clock), .in1(R11739));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11842 (.out1(R11843), .clock(clock), .in1(R11842));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11890 (.out1(R11891), .clock(clock), .in1(R11890));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11933 (.out1(R11934), .clock(clock), .in1(R11933));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12023 (.out1(R12024), .clock(clock), .in1(idx_3666));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1583 (.out1(_1532), .in1(R12024));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1584 (.out1(_1533), .in1(_1532), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3899 (.out1(R3900), .clock(clock), .in1(R3899));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4155 (.out1(R4156), .clock(clock), .in1(R4155));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4410 (.out1(R4411), .clock(clock), .in1(R4410));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4655 (.out1(R4656), .clock(clock), .in1(R4655));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4895 (.out1(R4896), .clock(clock), .in1(R4895));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5182 (.out1(R5183), .clock(clock), .in1(R5182));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5414 (.out1(R5415), .clock(clock), .in1(R5414));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5641 (.out1(R5642), .clock(clock), .in1(R5641));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5915 (.out1(R5916), .clock(clock), .in1(R5915));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6133 (.out1(R6134), .clock(clock), .in1(R6133));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6346 (.out1(R6347), .clock(clock), .in1(R6346));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6607 (.out1(R6608), .clock(clock), .in1(R6607));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6812 (.out1(R6813), .clock(clock), .in1(R6812));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7012 (.out1(R7013), .clock(clock), .in1(R7012));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7259 (.out1(R7260), .clock(clock), .in1(R7259));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7451 (.out1(R7452), .clock(clock), .in1(R7451));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7638 (.out1(R7639), .clock(clock), .in1(R7638));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7872 (.out1(R7873), .clock(clock), .in1(R7872));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8051 (.out1(R8052), .clock(clock), .in1(R8051));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8225 (.out1(R8226), .clock(clock), .in1(R8225));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8446 (.out1(R8447), .clock(clock), .in1(R8446));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8612 (.out1(R8613), .clock(clock), .in1(R8612));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8773 (.out1(R8774), .clock(clock), .in1(R8773));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8981 (.out1(R8982), .clock(clock), .in1(R8981));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9134 (.out1(R9135), .clock(clock), .in1(R9134));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9282 (.out1(R9283), .clock(clock), .in1(R9282));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9477 (.out1(R9478), .clock(clock), .in1(R9477));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9617 (.out1(R9618), .clock(clock), .in1(R9617));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9752 (.out1(R9753), .clock(clock), .in1(R9752));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9934 (.out1(R9935), .clock(clock), .in1(R9934));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10061 (.out1(R10062), .clock(clock), .in1(R10061));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10183 (.out1(R10184), .clock(clock), .in1(R10183));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10352 (.out1(R10353), .clock(clock), .in1(R10352));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10465 (.out1(R10466), .clock(clock), .in1(R10465));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10573 (.out1(R10574), .clock(clock), .in1(R10573));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10729 (.out1(R10730), .clock(clock), .in1(R10729));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10829 (.out1(R10830), .clock(clock), .in1(R10829));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10924 (.out1(R10925), .clock(clock), .in1(R10924));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11066 (.out1(R11067), .clock(clock), .in1(R11066));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11153 (.out1(R11154), .clock(clock), .in1(R11153));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11235 (.out1(R11236), .clock(clock), .in1(R11235));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11364 (.out1(R11365), .clock(clock), .in1(R11364));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11438 (.out1(R11439), .clock(clock), .in1(R11438));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11507 (.out1(R11508), .clock(clock), .in1(R11507));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11623 (.out1(R11624), .clock(clock), .in1(R11623));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11684 (.out1(R11685), .clock(clock), .in1(R11684));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11740 (.out1(R11741), .clock(clock), .in1(R11740));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11843 (.out1(R11844), .clock(clock), .in1(R11843));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11891 (.out1(R11892), .clock(clock), .in1(R11891));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11934 (.out1(R11935), .clock(clock), .in1(R11934));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12024 (.out1(R12025), .clock(clock), .in1(R12024));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12059 (.out1(R12060), .clock(clock), .in1(_1533));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1585 (.out1(_1534), .in1(vec112_3668_D), .in2(R12060));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3900 (.out1(R3901), .clock(clock), .in1(R3900));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4156 (.out1(R4157), .clock(clock), .in1(R4156));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4411 (.out1(R4412), .clock(clock), .in1(R4411));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4656 (.out1(R4657), .clock(clock), .in1(R4656));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4896 (.out1(R4897), .clock(clock), .in1(R4896));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5183 (.out1(R5184), .clock(clock), .in1(R5183));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5415 (.out1(R5416), .clock(clock), .in1(R5415));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5642 (.out1(R5643), .clock(clock), .in1(R5642));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5916 (.out1(R5917), .clock(clock), .in1(R5916));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6134 (.out1(R6135), .clock(clock), .in1(R6134));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6347 (.out1(R6348), .clock(clock), .in1(R6347));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6608 (.out1(R6609), .clock(clock), .in1(R6608));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6813 (.out1(R6814), .clock(clock), .in1(R6813));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7013 (.out1(R7014), .clock(clock), .in1(R7013));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7260 (.out1(R7261), .clock(clock), .in1(R7260));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7452 (.out1(R7453), .clock(clock), .in1(R7452));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7639 (.out1(R7640), .clock(clock), .in1(R7639));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7873 (.out1(R7874), .clock(clock), .in1(R7873));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8052 (.out1(R8053), .clock(clock), .in1(R8052));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8226 (.out1(R8227), .clock(clock), .in1(R8226));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8447 (.out1(R8448), .clock(clock), .in1(R8447));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8613 (.out1(R8614), .clock(clock), .in1(R8613));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8774 (.out1(R8775), .clock(clock), .in1(R8774));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8982 (.out1(R8983), .clock(clock), .in1(R8982));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9135 (.out1(R9136), .clock(clock), .in1(R9135));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9283 (.out1(R9284), .clock(clock), .in1(R9283));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9478 (.out1(R9479), .clock(clock), .in1(R9478));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9618 (.out1(R9619), .clock(clock), .in1(R9618));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9753 (.out1(R9754), .clock(clock), .in1(R9753));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9935 (.out1(R9936), .clock(clock), .in1(R9935));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10062 (.out1(R10063), .clock(clock), .in1(R10062));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10184 (.out1(R10185), .clock(clock), .in1(R10184));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10353 (.out1(R10354), .clock(clock), .in1(R10353));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10466 (.out1(R10467), .clock(clock), .in1(R10466));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10574 (.out1(R10575), .clock(clock), .in1(R10574));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10730 (.out1(R10731), .clock(clock), .in1(R10730));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10830 (.out1(R10831), .clock(clock), .in1(R10830));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10925 (.out1(R10926), .clock(clock), .in1(R10925));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11067 (.out1(R11068), .clock(clock), .in1(R11067));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11154 (.out1(R11155), .clock(clock), .in1(R11154));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11236 (.out1(R11237), .clock(clock), .in1(R11236));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11365 (.out1(R11366), .clock(clock), .in1(R11365));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11439 (.out1(R11440), .clock(clock), .in1(R11439));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11508 (.out1(R11509), .clock(clock), .in1(R11508));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11624 (.out1(R11625), .clock(clock), .in1(R11624));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11685 (.out1(R11686), .clock(clock), .in1(R11685));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11741 (.out1(R11742), .clock(clock), .in1(R11741));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11844 (.out1(R11845), .clock(clock), .in1(R11844));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11892 (.out1(R11893), .clock(clock), .in1(R11892));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11935 (.out1(R11936), .clock(clock), .in1(R11935));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12025 (.out1(R12026), .clock(clock), .in1(R12025));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12060 (.out1(R12061), .clock(clock), .in1(_1534));
  SRAM op1586 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1535),.ADR(R12061));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3901 (.out1(R3902), .clock(clock), .in1(R3901));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4157 (.out1(R4158), .clock(clock), .in1(R4157));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4412 (.out1(R4413), .clock(clock), .in1(R4412));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4657 (.out1(R4658), .clock(clock), .in1(R4657));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4897 (.out1(R4898), .clock(clock), .in1(R4897));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5184 (.out1(R5185), .clock(clock), .in1(R5184));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5416 (.out1(R5417), .clock(clock), .in1(R5416));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5643 (.out1(R5644), .clock(clock), .in1(R5643));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5917 (.out1(R5918), .clock(clock), .in1(R5917));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6135 (.out1(R6136), .clock(clock), .in1(R6135));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6348 (.out1(R6349), .clock(clock), .in1(R6348));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6609 (.out1(R6610), .clock(clock), .in1(R6609));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6814 (.out1(R6815), .clock(clock), .in1(R6814));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7014 (.out1(R7015), .clock(clock), .in1(R7014));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7261 (.out1(R7262), .clock(clock), .in1(R7261));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7453 (.out1(R7454), .clock(clock), .in1(R7453));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7640 (.out1(R7641), .clock(clock), .in1(R7640));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7874 (.out1(R7875), .clock(clock), .in1(R7874));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8053 (.out1(R8054), .clock(clock), .in1(R8053));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8227 (.out1(R8228), .clock(clock), .in1(R8227));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8448 (.out1(R8449), .clock(clock), .in1(R8448));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8614 (.out1(R8615), .clock(clock), .in1(R8614));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8775 (.out1(R8776), .clock(clock), .in1(R8775));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8983 (.out1(R8984), .clock(clock), .in1(R8983));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9136 (.out1(R9137), .clock(clock), .in1(R9136));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9284 (.out1(R9285), .clock(clock), .in1(R9284));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9479 (.out1(R9480), .clock(clock), .in1(R9479));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9619 (.out1(R9620), .clock(clock), .in1(R9619));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9754 (.out1(R9755), .clock(clock), .in1(R9754));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9936 (.out1(R9937), .clock(clock), .in1(R9936));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10063 (.out1(R10064), .clock(clock), .in1(R10063));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10185 (.out1(R10186), .clock(clock), .in1(R10185));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10354 (.out1(R10355), .clock(clock), .in1(R10354));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10467 (.out1(R10468), .clock(clock), .in1(R10467));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10575 (.out1(R10576), .clock(clock), .in1(R10575));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10731 (.out1(R10732), .clock(clock), .in1(R10731));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10831 (.out1(R10832), .clock(clock), .in1(R10831));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10926 (.out1(R10927), .clock(clock), .in1(R10926));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11068 (.out1(R11069), .clock(clock), .in1(R11068));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11155 (.out1(R11156), .clock(clock), .in1(R11155));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11237 (.out1(R11238), .clock(clock), .in1(R11237));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11366 (.out1(R11367), .clock(clock), .in1(R11366));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11440 (.out1(R11441), .clock(clock), .in1(R11440));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11509 (.out1(R11510), .clock(clock), .in1(R11509));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11625 (.out1(R11626), .clock(clock), .in1(R11625));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11686 (.out1(R11687), .clock(clock), .in1(R11686));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11742 (.out1(R11743), .clock(clock), .in1(R11742));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11845 (.out1(R11846), .clock(clock), .in1(R11845));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11893 (.out1(R11894), .clock(clock), .in1(R11893));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11936 (.out1(R11937), .clock(clock), .in1(R11936));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12026 (.out1(R12027), .clock(clock), .in1(R12026));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12061 (.out1(R12062), .clock(clock), .in1(_1535));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(4), .BITSIZE_out1(64), .PRECISION(64)) op1580 (.out1(_1530), .in1(ip2_3602_D), .in2(4 'd 10));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1581 (.out1(_1531), .in1(_1530));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op1582 (.out1(off_3667), .in1(_1531), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1587 (.out1(_1536), .in1(R12062), .in2(off_3667));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3902 (.out1(R3903), .clock(clock), .in1(R3902));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4158 (.out1(R4159), .clock(clock), .in1(R4158));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4413 (.out1(R4414), .clock(clock), .in1(R4413));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4658 (.out1(R4659), .clock(clock), .in1(R4658));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4898 (.out1(R4899), .clock(clock), .in1(R4898));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5185 (.out1(R5186), .clock(clock), .in1(R5185));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5417 (.out1(R5418), .clock(clock), .in1(R5417));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5644 (.out1(R5645), .clock(clock), .in1(R5644));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5918 (.out1(R5919), .clock(clock), .in1(R5918));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6136 (.out1(R6137), .clock(clock), .in1(R6136));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6349 (.out1(R6350), .clock(clock), .in1(R6349));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6610 (.out1(R6611), .clock(clock), .in1(R6610));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6815 (.out1(R6816), .clock(clock), .in1(R6815));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7015 (.out1(R7016), .clock(clock), .in1(R7015));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7262 (.out1(R7263), .clock(clock), .in1(R7262));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7454 (.out1(R7455), .clock(clock), .in1(R7454));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7641 (.out1(R7642), .clock(clock), .in1(R7641));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7875 (.out1(R7876), .clock(clock), .in1(R7875));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8054 (.out1(R8055), .clock(clock), .in1(R8054));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8228 (.out1(R8229), .clock(clock), .in1(R8228));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8449 (.out1(R8450), .clock(clock), .in1(R8449));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8615 (.out1(R8616), .clock(clock), .in1(R8615));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8776 (.out1(R8777), .clock(clock), .in1(R8776));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8984 (.out1(R8985), .clock(clock), .in1(R8984));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9137 (.out1(R9138), .clock(clock), .in1(R9137));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9285 (.out1(R9286), .clock(clock), .in1(R9285));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9480 (.out1(R9481), .clock(clock), .in1(R9480));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9620 (.out1(R9621), .clock(clock), .in1(R9620));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9755 (.out1(R9756), .clock(clock), .in1(R9755));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9937 (.out1(R9938), .clock(clock), .in1(R9937));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10064 (.out1(R10065), .clock(clock), .in1(R10064));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10186 (.out1(R10187), .clock(clock), .in1(R10186));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10355 (.out1(R10356), .clock(clock), .in1(R10355));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10468 (.out1(R10469), .clock(clock), .in1(R10468));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10576 (.out1(R10577), .clock(clock), .in1(R10576));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10732 (.out1(R10733), .clock(clock), .in1(R10732));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10832 (.out1(R10833), .clock(clock), .in1(R10832));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10927 (.out1(R10928), .clock(clock), .in1(R10927));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11069 (.out1(R11070), .clock(clock), .in1(R11069));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11156 (.out1(R11157), .clock(clock), .in1(R11156));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11238 (.out1(R11239), .clock(clock), .in1(R11238));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11367 (.out1(R11368), .clock(clock), .in1(R11367));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11441 (.out1(R11442), .clock(clock), .in1(R11441));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11510 (.out1(R11511), .clock(clock), .in1(R11510));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11626 (.out1(R11627), .clock(clock), .in1(R11626));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11687 (.out1(R11688), .clock(clock), .in1(R11687));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11743 (.out1(R11744), .clock(clock), .in1(R11743));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11846 (.out1(R11847), .clock(clock), .in1(R11846));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11894 (.out1(R11895), .clock(clock), .in1(R11894));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11937 (.out1(R11938), .clock(clock), .in1(R11937));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12027 (.out1(R12028), .clock(clock), .in1(R12027));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12062 (.out1(R12063), .clock(clock), .in1(off_3667));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12092 (.out1(R12093), .clock(clock), .in1(_1536));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op1588 (.out1(_1537), .in1(R12093), .in2(1 'd 1));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op1589 (.out1(ifout1589), .in1(_1537), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1657 (.out1(_1605), .in1(R12028));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1650 (.out1(_1598), .in1(R12028));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1639 (.out1(_1587), .in1(R12028));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1619 (.out1(_1567), .in1(R12028));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1658 (.out1(_1606), .in1(_1605), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1651 (.out1(_1599), .in1(_1598), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1640 (.out1(_1588), .in1(_1587), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1620 (.out1(_1568), .in1(_1567), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3903 (.out1(R3904), .clock(clock), .in1(R3903));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4159 (.out1(R4160), .clock(clock), .in1(R4159));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4414 (.out1(R4415), .clock(clock), .in1(R4414));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4659 (.out1(R4660), .clock(clock), .in1(R4659));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4899 (.out1(R4900), .clock(clock), .in1(R4899));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5186 (.out1(R5187), .clock(clock), .in1(R5186));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5418 (.out1(R5419), .clock(clock), .in1(R5418));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5645 (.out1(R5646), .clock(clock), .in1(R5645));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5919 (.out1(R5920), .clock(clock), .in1(R5919));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6137 (.out1(R6138), .clock(clock), .in1(R6137));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6350 (.out1(R6351), .clock(clock), .in1(R6350));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6611 (.out1(R6612), .clock(clock), .in1(R6611));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6816 (.out1(R6817), .clock(clock), .in1(R6816));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7016 (.out1(R7017), .clock(clock), .in1(R7016));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7263 (.out1(R7264), .clock(clock), .in1(R7263));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7455 (.out1(R7456), .clock(clock), .in1(R7455));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7642 (.out1(R7643), .clock(clock), .in1(R7642));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7876 (.out1(R7877), .clock(clock), .in1(R7876));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8055 (.out1(R8056), .clock(clock), .in1(R8055));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8229 (.out1(R8230), .clock(clock), .in1(R8229));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8450 (.out1(R8451), .clock(clock), .in1(R8450));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8616 (.out1(R8617), .clock(clock), .in1(R8616));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8777 (.out1(R8778), .clock(clock), .in1(R8777));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8985 (.out1(R8986), .clock(clock), .in1(R8985));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9138 (.out1(R9139), .clock(clock), .in1(R9138));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9286 (.out1(R9287), .clock(clock), .in1(R9286));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9481 (.out1(R9482), .clock(clock), .in1(R9481));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9621 (.out1(R9622), .clock(clock), .in1(R9621));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9756 (.out1(R9757), .clock(clock), .in1(R9756));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9938 (.out1(R9939), .clock(clock), .in1(R9938));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10065 (.out1(R10066), .clock(clock), .in1(R10065));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10187 (.out1(R10188), .clock(clock), .in1(R10187));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10356 (.out1(R10357), .clock(clock), .in1(R10356));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10469 (.out1(R10470), .clock(clock), .in1(R10469));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10577 (.out1(R10578), .clock(clock), .in1(R10577));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10733 (.out1(R10734), .clock(clock), .in1(R10733));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10833 (.out1(R10834), .clock(clock), .in1(R10833));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10928 (.out1(R10929), .clock(clock), .in1(R10928));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11070 (.out1(R11071), .clock(clock), .in1(R11070));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11157 (.out1(R11158), .clock(clock), .in1(R11157));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11239 (.out1(R11240), .clock(clock), .in1(R11239));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11368 (.out1(R11369), .clock(clock), .in1(R11368));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11442 (.out1(R11443), .clock(clock), .in1(R11442));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11511 (.out1(R11512), .clock(clock), .in1(R11511));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11627 (.out1(R11628), .clock(clock), .in1(R11627));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11688 (.out1(R11689), .clock(clock), .in1(R11688));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11744 (.out1(R11745), .clock(clock), .in1(R11744));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11847 (.out1(R11848), .clock(clock), .in1(R11847));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11895 (.out1(R11896), .clock(clock), .in1(R11895));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11938 (.out1(R11939), .clock(clock), .in1(R11938));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12028 (.out1(R12029), .clock(clock), .in1(R12028));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12063 (.out1(R12064), .clock(clock), .in1(R12063));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12093 (.out1(R12094), .clock(clock), .in1(ifout1589));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12130 (.out1(R12131), .clock(clock), .in1(_1606));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12131 (.out1(R12132), .clock(clock), .in1(_1599));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12132 (.out1(R12133), .clock(clock), .in1(_1588));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12133 (.out1(R12134), .clock(clock), .in1(_1568));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1632 (.out1(_1580), .in1(R12029));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1612 (.out1(_1560), .in1(R12029));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1601 (.out1(_1549), .in1(R12029));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1594 (.out1(_1542), .in1(R12029));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1661 (.out1(_1609), .in1(2 'd 2), .in2(R12064));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1633 (.out1(_1581), .in1(_1580), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1613 (.out1(_1561), .in1(_1560), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1602 (.out1(_1550), .in1(_1549), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1595 (.out1(_1543), .in1(_1542), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1659 (.out1(_1607), .in1(vec112_3668_D), .in2(R12131));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1652 (.out1(_1600), .in1(vec112_3668_D), .in2(R12132));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1641 (.out1(_1589), .in1(vec112_3668_D), .in2(R12133));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1621 (.out1(_1569), .in1(vec112_3668_D), .in2(R12134));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3904 (.out1(R3905), .clock(clock), .in1(R3904));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4160 (.out1(R4161), .clock(clock), .in1(R4160));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4415 (.out1(R4416), .clock(clock), .in1(R4415));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4660 (.out1(R4661), .clock(clock), .in1(R4660));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4900 (.out1(R4901), .clock(clock), .in1(R4900));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5187 (.out1(R5188), .clock(clock), .in1(R5187));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5419 (.out1(R5420), .clock(clock), .in1(R5419));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5646 (.out1(R5647), .clock(clock), .in1(R5646));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5920 (.out1(R5921), .clock(clock), .in1(R5920));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6138 (.out1(R6139), .clock(clock), .in1(R6138));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6351 (.out1(R6352), .clock(clock), .in1(R6351));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6612 (.out1(R6613), .clock(clock), .in1(R6612));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6817 (.out1(R6818), .clock(clock), .in1(R6817));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7017 (.out1(R7018), .clock(clock), .in1(R7017));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7264 (.out1(R7265), .clock(clock), .in1(R7264));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7456 (.out1(R7457), .clock(clock), .in1(R7456));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7643 (.out1(R7644), .clock(clock), .in1(R7643));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7877 (.out1(R7878), .clock(clock), .in1(R7877));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8056 (.out1(R8057), .clock(clock), .in1(R8056));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8230 (.out1(R8231), .clock(clock), .in1(R8230));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8451 (.out1(R8452), .clock(clock), .in1(R8451));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8617 (.out1(R8618), .clock(clock), .in1(R8617));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8778 (.out1(R8779), .clock(clock), .in1(R8778));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8986 (.out1(R8987), .clock(clock), .in1(R8986));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9139 (.out1(R9140), .clock(clock), .in1(R9139));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9287 (.out1(R9288), .clock(clock), .in1(R9287));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9482 (.out1(R9483), .clock(clock), .in1(R9482));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9622 (.out1(R9623), .clock(clock), .in1(R9622));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9757 (.out1(R9758), .clock(clock), .in1(R9757));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9939 (.out1(R9940), .clock(clock), .in1(R9939));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10066 (.out1(R10067), .clock(clock), .in1(R10066));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10188 (.out1(R10189), .clock(clock), .in1(R10188));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10357 (.out1(R10358), .clock(clock), .in1(R10357));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10470 (.out1(R10471), .clock(clock), .in1(R10470));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10578 (.out1(R10579), .clock(clock), .in1(R10578));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10734 (.out1(R10735), .clock(clock), .in1(R10734));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10834 (.out1(R10835), .clock(clock), .in1(R10834));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10929 (.out1(R10930), .clock(clock), .in1(R10929));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11071 (.out1(R11072), .clock(clock), .in1(R11071));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11158 (.out1(R11159), .clock(clock), .in1(R11158));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11240 (.out1(R11241), .clock(clock), .in1(R11240));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11369 (.out1(R11370), .clock(clock), .in1(R11369));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11443 (.out1(R11444), .clock(clock), .in1(R11443));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11512 (.out1(R11513), .clock(clock), .in1(R11512));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11628 (.out1(R11629), .clock(clock), .in1(R11628));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11689 (.out1(R11690), .clock(clock), .in1(R11689));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11745 (.out1(R11746), .clock(clock), .in1(R11745));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11848 (.out1(R11849), .clock(clock), .in1(R11848));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11896 (.out1(R11897), .clock(clock), .in1(R11896));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11939 (.out1(R11940), .clock(clock), .in1(R11939));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12029 (.out1(R12030), .clock(clock), .in1(R12029));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12064 (.out1(R12065), .clock(clock), .in1(R12064));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12094 (.out1(R12095), .clock(clock), .in1(R12094));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12134 (.out1(R12135), .clock(clock), .in1(_1609));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12135 (.out1(R12136), .clock(clock), .in1(_1581));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12136 (.out1(R12137), .clock(clock), .in1(_1561));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12137 (.out1(R12138), .clock(clock), .in1(_1550));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12138 (.out1(R12139), .clock(clock), .in1(_1543));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12139 (.out1(R12140), .clock(clock), .in1(_1607));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12140 (.out1(R12141), .clock(clock), .in1(_1600));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12141 (.out1(R12142), .clock(clock), .in1(_1589));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12142 (.out1(R12143), .clock(clock), .in1(_1569));
  SRAM op1660 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1608),.ADR(R12140));
  SRAM op1653 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1601),.ADR(R12141));
  SRAM op1642 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1590),.ADR(R12142));
  SRAM op1622 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1570),.ADR(R12143));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1654 (.out1(_1602), .in1(2 'd 2), .in2(R12065));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1643 (.out1(_1591), .in1(2 'd 2), .in2(R12065));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1636 (.out1(_1584), .in1(2 'd 2), .in2(R12065));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1623 (.out1(_1571), .in1(2 'd 2), .in2(R12065));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1616 (.out1(_1564), .in1(2 'd 2), .in2(R12065));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1605 (.out1(_1553), .in1(2 'd 2), .in2(R12065));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1634 (.out1(_1582), .in1(vec112_3668_D), .in2(R12136));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1614 (.out1(_1562), .in1(vec112_3668_D), .in2(R12137));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1603 (.out1(_1551), .in1(vec112_3668_D), .in2(R12138));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1596 (.out1(_1544), .in1(vec112_3668_D), .in2(R12139));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1662 (.out1(_1610), .in1(R12135), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3905 (.out1(R3906), .clock(clock), .in1(R3905));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4161 (.out1(R4162), .clock(clock), .in1(R4161));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4416 (.out1(R4417), .clock(clock), .in1(R4416));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4661 (.out1(R4662), .clock(clock), .in1(R4661));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4901 (.out1(R4902), .clock(clock), .in1(R4901));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5188 (.out1(R5189), .clock(clock), .in1(R5188));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5420 (.out1(R5421), .clock(clock), .in1(R5420));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5647 (.out1(R5648), .clock(clock), .in1(R5647));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5921 (.out1(R5922), .clock(clock), .in1(R5921));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6139 (.out1(R6140), .clock(clock), .in1(R6139));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6352 (.out1(R6353), .clock(clock), .in1(R6352));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6613 (.out1(R6614), .clock(clock), .in1(R6613));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6818 (.out1(R6819), .clock(clock), .in1(R6818));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7018 (.out1(R7019), .clock(clock), .in1(R7018));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7265 (.out1(R7266), .clock(clock), .in1(R7265));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7457 (.out1(R7458), .clock(clock), .in1(R7457));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7644 (.out1(R7645), .clock(clock), .in1(R7644));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7878 (.out1(R7879), .clock(clock), .in1(R7878));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8057 (.out1(R8058), .clock(clock), .in1(R8057));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8231 (.out1(R8232), .clock(clock), .in1(R8231));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8452 (.out1(R8453), .clock(clock), .in1(R8452));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8618 (.out1(R8619), .clock(clock), .in1(R8618));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8779 (.out1(R8780), .clock(clock), .in1(R8779));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8987 (.out1(R8988), .clock(clock), .in1(R8987));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9140 (.out1(R9141), .clock(clock), .in1(R9140));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9288 (.out1(R9289), .clock(clock), .in1(R9288));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9483 (.out1(R9484), .clock(clock), .in1(R9483));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9623 (.out1(R9624), .clock(clock), .in1(R9623));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9758 (.out1(R9759), .clock(clock), .in1(R9758));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9940 (.out1(R9941), .clock(clock), .in1(R9940));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10067 (.out1(R10068), .clock(clock), .in1(R10067));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10189 (.out1(R10190), .clock(clock), .in1(R10189));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10358 (.out1(R10359), .clock(clock), .in1(R10358));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10471 (.out1(R10472), .clock(clock), .in1(R10471));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10579 (.out1(R10580), .clock(clock), .in1(R10579));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10735 (.out1(R10736), .clock(clock), .in1(R10735));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10835 (.out1(R10836), .clock(clock), .in1(R10835));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10930 (.out1(R10931), .clock(clock), .in1(R10930));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11072 (.out1(R11073), .clock(clock), .in1(R11072));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11159 (.out1(R11160), .clock(clock), .in1(R11159));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11241 (.out1(R11242), .clock(clock), .in1(R11241));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11370 (.out1(R11371), .clock(clock), .in1(R11370));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11444 (.out1(R11445), .clock(clock), .in1(R11444));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11513 (.out1(R11514), .clock(clock), .in1(R11513));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11629 (.out1(R11630), .clock(clock), .in1(R11629));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11690 (.out1(R11691), .clock(clock), .in1(R11690));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11746 (.out1(R11747), .clock(clock), .in1(R11746));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11849 (.out1(R11850), .clock(clock), .in1(R11849));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11897 (.out1(R11898), .clock(clock), .in1(R11897));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11940 (.out1(R11941), .clock(clock), .in1(R11940));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12030 (.out1(R12031), .clock(clock), .in1(R12030));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12065 (.out1(R12066), .clock(clock), .in1(R12065));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12095 (.out1(R12096), .clock(clock), .in1(R12095));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12143 (.out1(R12144), .clock(clock), .in1(_1608));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12144 (.out1(R12145), .clock(clock), .in1(_1601));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12145 (.out1(R12146), .clock(clock), .in1(_1590));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12146 (.out1(R12147), .clock(clock), .in1(_1570));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12147 (.out1(R12148), .clock(clock), .in1(_1602));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12148 (.out1(R12149), .clock(clock), .in1(_1591));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12149 (.out1(R12150), .clock(clock), .in1(_1584));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12150 (.out1(R12151), .clock(clock), .in1(_1571));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12151 (.out1(R12152), .clock(clock), .in1(_1564));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12152 (.out1(R12153), .clock(clock), .in1(_1553));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12153 (.out1(R12154), .clock(clock), .in1(_1582));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12154 (.out1(R12155), .clock(clock), .in1(_1562));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12155 (.out1(R12156), .clock(clock), .in1(_1551));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12156 (.out1(R12157), .clock(clock), .in1(_1544));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12157 (.out1(R12158), .clock(clock), .in1(_1610));
  SRAM op1635 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1583),.ADR(R12154));
  SRAM op1615 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1563),.ADR(R12155));
  SRAM op1604 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1552),.ADR(R12156));
  SRAM op1597 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1545),.ADR(R12157));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1663 (.out1(_1611), .in1(R12144), .in2(R12158));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1664 (.out1(_1612), .in1(_1611), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1655 (.out1(_1603), .in1(R12148), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1644 (.out1(_1592), .in1(R12149), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1624 (.out1(_1572), .in1(R12151), .in2(64 'd 18446744073709551615));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1598 (.out1(_1546), .in1(2 'd 2), .in2(R12066));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1665 (.out1(_1613), .in1(_1612), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1656 (.out1(_1604), .in1(R12145), .in2(_1603));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1645 (.out1(_1593), .in1(R12146), .in2(_1592));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1625 (.out1(_1573), .in1(R12147), .in2(_1572));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1666 (.out1(_1614), .in1(_1604), .in2(_1613));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1646 (.out1(_1594), .in1(_1593), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1637 (.out1(_1585), .in1(R12150), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1626 (.out1(_1574), .in1(_1573), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1617 (.out1(_1565), .in1(R12152), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1606 (.out1(_1554), .in1(R12153), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3906 (.out1(R3907), .clock(clock), .in1(R3906));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4162 (.out1(R4163), .clock(clock), .in1(R4162));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4417 (.out1(R4418), .clock(clock), .in1(R4417));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4662 (.out1(R4663), .clock(clock), .in1(R4662));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4902 (.out1(R4903), .clock(clock), .in1(R4902));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5189 (.out1(R5190), .clock(clock), .in1(R5189));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5421 (.out1(R5422), .clock(clock), .in1(R5421));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5648 (.out1(R5649), .clock(clock), .in1(R5648));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5922 (.out1(R5923), .clock(clock), .in1(R5922));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6140 (.out1(R6141), .clock(clock), .in1(R6140));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6353 (.out1(R6354), .clock(clock), .in1(R6353));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6614 (.out1(R6615), .clock(clock), .in1(R6614));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6819 (.out1(R6820), .clock(clock), .in1(R6819));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7019 (.out1(R7020), .clock(clock), .in1(R7019));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7266 (.out1(R7267), .clock(clock), .in1(R7266));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7458 (.out1(R7459), .clock(clock), .in1(R7458));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7645 (.out1(R7646), .clock(clock), .in1(R7645));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7879 (.out1(R7880), .clock(clock), .in1(R7879));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8058 (.out1(R8059), .clock(clock), .in1(R8058));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8232 (.out1(R8233), .clock(clock), .in1(R8232));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8453 (.out1(R8454), .clock(clock), .in1(R8453));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8619 (.out1(R8620), .clock(clock), .in1(R8619));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8780 (.out1(R8781), .clock(clock), .in1(R8780));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8988 (.out1(R8989), .clock(clock), .in1(R8988));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9141 (.out1(R9142), .clock(clock), .in1(R9141));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9289 (.out1(R9290), .clock(clock), .in1(R9289));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9484 (.out1(R9485), .clock(clock), .in1(R9484));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9624 (.out1(R9625), .clock(clock), .in1(R9624));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9759 (.out1(R9760), .clock(clock), .in1(R9759));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9941 (.out1(R9942), .clock(clock), .in1(R9941));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10068 (.out1(R10069), .clock(clock), .in1(R10068));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10190 (.out1(R10191), .clock(clock), .in1(R10190));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10359 (.out1(R10360), .clock(clock), .in1(R10359));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10472 (.out1(R10473), .clock(clock), .in1(R10472));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10580 (.out1(R10581), .clock(clock), .in1(R10580));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10736 (.out1(R10737), .clock(clock), .in1(R10736));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10836 (.out1(R10837), .clock(clock), .in1(R10836));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10931 (.out1(R10932), .clock(clock), .in1(R10931));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11073 (.out1(R11074), .clock(clock), .in1(R11073));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11160 (.out1(R11161), .clock(clock), .in1(R11160));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11242 (.out1(R11243), .clock(clock), .in1(R11242));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11371 (.out1(R11372), .clock(clock), .in1(R11371));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11445 (.out1(R11446), .clock(clock), .in1(R11445));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11514 (.out1(R11515), .clock(clock), .in1(R11514));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11630 (.out1(R11631), .clock(clock), .in1(R11630));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11691 (.out1(R11692), .clock(clock), .in1(R11691));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11747 (.out1(R11748), .clock(clock), .in1(R11747));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11850 (.out1(R11851), .clock(clock), .in1(R11850));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11898 (.out1(R11899), .clock(clock), .in1(R11898));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11941 (.out1(R11942), .clock(clock), .in1(R11941));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12031 (.out1(R12032), .clock(clock), .in1(R12031));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12066 (.out1(R12067), .clock(clock), .in1(R12066));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12096 (.out1(R12097), .clock(clock), .in1(R12096));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12158 (.out1(R12159), .clock(clock), .in1(_1583));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12159 (.out1(R12160), .clock(clock), .in1(_1563));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12160 (.out1(R12161), .clock(clock), .in1(_1552));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12161 (.out1(R12162), .clock(clock), .in1(_1545));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12162 (.out1(R12163), .clock(clock), .in1(_1546));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12163 (.out1(R12164), .clock(clock), .in1(_1614));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12164 (.out1(R12165), .clock(clock), .in1(_1594));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12165 (.out1(R12166), .clock(clock), .in1(_1585));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12166 (.out1(R12167), .clock(clock), .in1(_1574));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12167 (.out1(R12168), .clock(clock), .in1(_1565));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12168 (.out1(R12169), .clock(clock), .in1(_1554));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1647 (.out1(_1595), .in1(R12165), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1638 (.out1(_1586), .in1(R12159), .in2(R12166));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1607 (.out1(_1555), .in1(R12161), .in2(R12169));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1667 (.out1(_1615), .in1(R12164), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1648 (.out1(_1596), .in1(_1586), .in2(_1595));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1627 (.out1(_1575), .in1(R12167), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1618 (.out1(_1566), .in1(R12160), .in2(R12168));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1608 (.out1(_1556), .in1(_1555), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1599 (.out1(_1547), .in1(R12163), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1628 (.out1(_1576), .in1(_1566), .in2(_1575));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1668 (.out1(_1616), .in1(_1615), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1649 (.out1(_1597), .in1(_1596), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1609 (.out1(_1557), .in1(_1556), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1600 (.out1(_1548), .in1(R12162), .in2(_1547));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1669 (.out1(_1617), .in1(_1597), .in2(_1616));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1629 (.out1(_1577), .in1(_1576), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1610 (.out1(_1558), .in1(_1548), .in2(_1557));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3907 (.out1(R3908), .clock(clock), .in1(R3907));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4163 (.out1(R4164), .clock(clock), .in1(R4163));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4418 (.out1(R4419), .clock(clock), .in1(R4418));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4663 (.out1(R4664), .clock(clock), .in1(R4663));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4903 (.out1(R4904), .clock(clock), .in1(R4903));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5190 (.out1(R5191), .clock(clock), .in1(R5190));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5422 (.out1(R5423), .clock(clock), .in1(R5422));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5649 (.out1(R5650), .clock(clock), .in1(R5649));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5923 (.out1(R5924), .clock(clock), .in1(R5923));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6141 (.out1(R6142), .clock(clock), .in1(R6141));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6354 (.out1(R6355), .clock(clock), .in1(R6354));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6615 (.out1(R6616), .clock(clock), .in1(R6615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6820 (.out1(R6821), .clock(clock), .in1(R6820));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7020 (.out1(R7021), .clock(clock), .in1(R7020));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7267 (.out1(R7268), .clock(clock), .in1(R7267));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7459 (.out1(R7460), .clock(clock), .in1(R7459));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7646 (.out1(R7647), .clock(clock), .in1(R7646));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7880 (.out1(R7881), .clock(clock), .in1(R7880));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8059 (.out1(R8060), .clock(clock), .in1(R8059));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8233 (.out1(R8234), .clock(clock), .in1(R8233));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8454 (.out1(R8455), .clock(clock), .in1(R8454));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8620 (.out1(R8621), .clock(clock), .in1(R8620));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8781 (.out1(R8782), .clock(clock), .in1(R8781));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8989 (.out1(R8990), .clock(clock), .in1(R8989));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9142 (.out1(R9143), .clock(clock), .in1(R9142));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9290 (.out1(R9291), .clock(clock), .in1(R9290));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9485 (.out1(R9486), .clock(clock), .in1(R9485));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9625 (.out1(R9626), .clock(clock), .in1(R9625));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9760 (.out1(R9761), .clock(clock), .in1(R9760));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9942 (.out1(R9943), .clock(clock), .in1(R9942));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10069 (.out1(R10070), .clock(clock), .in1(R10069));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10191 (.out1(R10192), .clock(clock), .in1(R10191));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10360 (.out1(R10361), .clock(clock), .in1(R10360));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10473 (.out1(R10474), .clock(clock), .in1(R10473));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10581 (.out1(R10582), .clock(clock), .in1(R10581));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10737 (.out1(R10738), .clock(clock), .in1(R10737));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10837 (.out1(R10838), .clock(clock), .in1(R10837));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10932 (.out1(R10933), .clock(clock), .in1(R10932));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11074 (.out1(R11075), .clock(clock), .in1(R11074));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11161 (.out1(R11162), .clock(clock), .in1(R11161));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11243 (.out1(R11244), .clock(clock), .in1(R11243));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11372 (.out1(R11373), .clock(clock), .in1(R11372));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11446 (.out1(R11447), .clock(clock), .in1(R11446));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11515 (.out1(R11516), .clock(clock), .in1(R11515));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11631 (.out1(R11632), .clock(clock), .in1(R11631));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11692 (.out1(R11693), .clock(clock), .in1(R11692));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11748 (.out1(R11749), .clock(clock), .in1(R11748));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11851 (.out1(R11852), .clock(clock), .in1(R11851));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11899 (.out1(R11900), .clock(clock), .in1(R11899));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11942 (.out1(R11943), .clock(clock), .in1(R11942));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12032 (.out1(R12033), .clock(clock), .in1(R12032));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12067 (.out1(R12068), .clock(clock), .in1(R12067));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12097 (.out1(R12098), .clock(clock), .in1(R12097));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12169 (.out1(R12170), .clock(clock), .in1(_1617));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12170 (.out1(R12171), .clock(clock), .in1(_1577));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12171 (.out1(R12172), .clock(clock), .in1(_1558));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1590 (.out1(_1538), .in1(R12033));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1630 (.out1(_1578), .in1(R12171), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1611 (.out1(_1559), .in1(R12172), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op1670 (.out1(_1618), .in1(R12170), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1631 (.out1(_1579), .in1(_1559), .in2(_1578));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1591 (.out1(_1539), .in1(_1538), .in2(2 'd 2));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1671 (.out1(_1619), .in1(_1579), .in2(_1618));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op1672 (.out1(_1620), .in1(_1619), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3908 (.out1(R3909), .clock(clock), .in1(R3908));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4164 (.out1(R4165), .clock(clock), .in1(R4164));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4419 (.out1(R4420), .clock(clock), .in1(R4419));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4664 (.out1(R4665), .clock(clock), .in1(R4664));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4904 (.out1(R4905), .clock(clock), .in1(R4904));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5191 (.out1(R5192), .clock(clock), .in1(R5191));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5423 (.out1(R5424), .clock(clock), .in1(R5423));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5650 (.out1(R5651), .clock(clock), .in1(R5650));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5924 (.out1(R5925), .clock(clock), .in1(R5924));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6142 (.out1(R6143), .clock(clock), .in1(R6142));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6355 (.out1(R6356), .clock(clock), .in1(R6355));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6616 (.out1(R6617), .clock(clock), .in1(R6616));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6821 (.out1(R6822), .clock(clock), .in1(R6821));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7021 (.out1(R7022), .clock(clock), .in1(R7021));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7268 (.out1(R7269), .clock(clock), .in1(R7268));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7460 (.out1(R7461), .clock(clock), .in1(R7460));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7647 (.out1(R7648), .clock(clock), .in1(R7647));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7881 (.out1(R7882), .clock(clock), .in1(R7881));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8060 (.out1(R8061), .clock(clock), .in1(R8060));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8234 (.out1(R8235), .clock(clock), .in1(R8234));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8455 (.out1(R8456), .clock(clock), .in1(R8455));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8621 (.out1(R8622), .clock(clock), .in1(R8621));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8782 (.out1(R8783), .clock(clock), .in1(R8782));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8990 (.out1(R8991), .clock(clock), .in1(R8990));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9143 (.out1(R9144), .clock(clock), .in1(R9143));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9291 (.out1(R9292), .clock(clock), .in1(R9291));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9486 (.out1(R9487), .clock(clock), .in1(R9486));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9626 (.out1(R9627), .clock(clock), .in1(R9626));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9761 (.out1(R9762), .clock(clock), .in1(R9761));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9943 (.out1(R9944), .clock(clock), .in1(R9943));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10070 (.out1(R10071), .clock(clock), .in1(R10070));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10192 (.out1(R10193), .clock(clock), .in1(R10192));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10361 (.out1(R10362), .clock(clock), .in1(R10361));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10474 (.out1(R10475), .clock(clock), .in1(R10474));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10582 (.out1(R10583), .clock(clock), .in1(R10582));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10738 (.out1(R10739), .clock(clock), .in1(R10738));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10838 (.out1(R10839), .clock(clock), .in1(R10838));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10933 (.out1(R10934), .clock(clock), .in1(R10933));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11075 (.out1(R11076), .clock(clock), .in1(R11075));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11162 (.out1(R11163), .clock(clock), .in1(R11162));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11244 (.out1(R11245), .clock(clock), .in1(R11244));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11373 (.out1(R11374), .clock(clock), .in1(R11373));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11447 (.out1(R11448), .clock(clock), .in1(R11447));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11516 (.out1(R11517), .clock(clock), .in1(R11516));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11632 (.out1(R11633), .clock(clock), .in1(R11632));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11693 (.out1(R11694), .clock(clock), .in1(R11693));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11749 (.out1(R11750), .clock(clock), .in1(R11749));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11852 (.out1(R11853), .clock(clock), .in1(R11852));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11900 (.out1(R11901), .clock(clock), .in1(R11900));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11943 (.out1(R11944), .clock(clock), .in1(R11943));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12033 (.out1(R12034), .clock(clock), .in1(R12033));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12068 (.out1(R12069), .clock(clock), .in1(R12068));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12098 (.out1(R12099), .clock(clock), .in1(R12098));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12172 (.out1(R12173), .clock(clock), .in1(_1539));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12173 (.out1(R12174), .clock(clock), .in1(_1620));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op1673 (.out1(_1621), .in1(R12174), .in2(57 'd 72340172838076673));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1592 (.out1(_1540), .in1(base0_112_3673_D), .in2(R12173));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3909 (.out1(R3910), .clock(clock), .in1(R3909));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4165 (.out1(R4166), .clock(clock), .in1(R4165));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4420 (.out1(R4421), .clock(clock), .in1(R4420));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4665 (.out1(R4666), .clock(clock), .in1(R4665));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4905 (.out1(R4906), .clock(clock), .in1(R4905));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5192 (.out1(R5193), .clock(clock), .in1(R5192));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5424 (.out1(R5425), .clock(clock), .in1(R5424));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5651 (.out1(R5652), .clock(clock), .in1(R5651));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5925 (.out1(R5926), .clock(clock), .in1(R5925));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6143 (.out1(R6144), .clock(clock), .in1(R6143));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6356 (.out1(R6357), .clock(clock), .in1(R6356));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6617 (.out1(R6618), .clock(clock), .in1(R6617));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6822 (.out1(R6823), .clock(clock), .in1(R6822));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7022 (.out1(R7023), .clock(clock), .in1(R7022));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7269 (.out1(R7270), .clock(clock), .in1(R7269));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7461 (.out1(R7462), .clock(clock), .in1(R7461));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7648 (.out1(R7649), .clock(clock), .in1(R7648));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7882 (.out1(R7883), .clock(clock), .in1(R7882));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8061 (.out1(R8062), .clock(clock), .in1(R8061));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8235 (.out1(R8236), .clock(clock), .in1(R8235));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8456 (.out1(R8457), .clock(clock), .in1(R8456));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8622 (.out1(R8623), .clock(clock), .in1(R8622));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8783 (.out1(R8784), .clock(clock), .in1(R8783));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8991 (.out1(R8992), .clock(clock), .in1(R8991));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9144 (.out1(R9145), .clock(clock), .in1(R9144));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9292 (.out1(R9293), .clock(clock), .in1(R9292));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9487 (.out1(R9488), .clock(clock), .in1(R9487));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9627 (.out1(R9628), .clock(clock), .in1(R9627));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9762 (.out1(R9763), .clock(clock), .in1(R9762));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9944 (.out1(R9945), .clock(clock), .in1(R9944));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10071 (.out1(R10072), .clock(clock), .in1(R10071));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10193 (.out1(R10194), .clock(clock), .in1(R10193));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10362 (.out1(R10363), .clock(clock), .in1(R10362));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10475 (.out1(R10476), .clock(clock), .in1(R10475));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10583 (.out1(R10584), .clock(clock), .in1(R10583));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10739 (.out1(R10740), .clock(clock), .in1(R10739));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10839 (.out1(R10840), .clock(clock), .in1(R10839));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10934 (.out1(R10935), .clock(clock), .in1(R10934));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11076 (.out1(R11077), .clock(clock), .in1(R11076));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11163 (.out1(R11164), .clock(clock), .in1(R11163));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11245 (.out1(R11246), .clock(clock), .in1(R11245));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11374 (.out1(R11375), .clock(clock), .in1(R11374));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11448 (.out1(R11449), .clock(clock), .in1(R11448));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11517 (.out1(R11518), .clock(clock), .in1(R11517));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11633 (.out1(R11634), .clock(clock), .in1(R11633));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11694 (.out1(R11695), .clock(clock), .in1(R11694));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11750 (.out1(R11751), .clock(clock), .in1(R11750));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11853 (.out1(R11854), .clock(clock), .in1(R11853));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11901 (.out1(R11902), .clock(clock), .in1(R11901));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11944 (.out1(R11945), .clock(clock), .in1(R11944));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12034 (.out1(R12035), .clock(clock), .in1(R12034));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12069 (.out1(R12070), .clock(clock), .in1(R12069));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12099 (.out1(R12100), .clock(clock), .in1(R12099));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12174 (.out1(R12175), .clock(clock), .in1(_1621));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12175 (.out1(R12176), .clock(clock), .in1(_1540));
  SRAM op1593 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1541),.ADR(R12176));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op1674 (.out1(_1622), .in1(R12175), .in2(6 'd 56));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3910 (.out1(R3911), .clock(clock), .in1(R3910));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4166 (.out1(R4167), .clock(clock), .in1(R4166));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4421 (.out1(R4422), .clock(clock), .in1(R4421));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4666 (.out1(R4667), .clock(clock), .in1(R4666));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4906 (.out1(R4907), .clock(clock), .in1(R4906));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5193 (.out1(R5194), .clock(clock), .in1(R5193));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5425 (.out1(R5426), .clock(clock), .in1(R5425));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5652 (.out1(R5653), .clock(clock), .in1(R5652));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5926 (.out1(R5927), .clock(clock), .in1(R5926));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6144 (.out1(R6145), .clock(clock), .in1(R6144));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6357 (.out1(R6358), .clock(clock), .in1(R6357));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6618 (.out1(R6619), .clock(clock), .in1(R6618));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6823 (.out1(R6824), .clock(clock), .in1(R6823));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7023 (.out1(R7024), .clock(clock), .in1(R7023));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7270 (.out1(R7271), .clock(clock), .in1(R7270));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7462 (.out1(R7463), .clock(clock), .in1(R7462));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7649 (.out1(R7650), .clock(clock), .in1(R7649));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7883 (.out1(R7884), .clock(clock), .in1(R7883));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8062 (.out1(R8063), .clock(clock), .in1(R8062));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8236 (.out1(R8237), .clock(clock), .in1(R8236));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8457 (.out1(R8458), .clock(clock), .in1(R8457));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8623 (.out1(R8624), .clock(clock), .in1(R8623));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8784 (.out1(R8785), .clock(clock), .in1(R8784));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8992 (.out1(R8993), .clock(clock), .in1(R8992));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9145 (.out1(R9146), .clock(clock), .in1(R9145));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9293 (.out1(R9294), .clock(clock), .in1(R9293));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9488 (.out1(R9489), .clock(clock), .in1(R9488));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9628 (.out1(R9629), .clock(clock), .in1(R9628));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9763 (.out1(R9764), .clock(clock), .in1(R9763));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9945 (.out1(R9946), .clock(clock), .in1(R9945));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10072 (.out1(R10073), .clock(clock), .in1(R10072));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10194 (.out1(R10195), .clock(clock), .in1(R10194));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10363 (.out1(R10364), .clock(clock), .in1(R10363));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10476 (.out1(R10477), .clock(clock), .in1(R10476));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10584 (.out1(R10585), .clock(clock), .in1(R10584));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10740 (.out1(R10741), .clock(clock), .in1(R10740));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10840 (.out1(R10841), .clock(clock), .in1(R10840));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10935 (.out1(R10936), .clock(clock), .in1(R10935));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11077 (.out1(R11078), .clock(clock), .in1(R11077));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11164 (.out1(R11165), .clock(clock), .in1(R11164));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11246 (.out1(R11247), .clock(clock), .in1(R11246));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11375 (.out1(R11376), .clock(clock), .in1(R11375));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11449 (.out1(R11450), .clock(clock), .in1(R11449));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11518 (.out1(R11519), .clock(clock), .in1(R11518));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11634 (.out1(R11635), .clock(clock), .in1(R11634));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11695 (.out1(R11696), .clock(clock), .in1(R11695));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11751 (.out1(R11752), .clock(clock), .in1(R11751));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11854 (.out1(R11855), .clock(clock), .in1(R11854));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11902 (.out1(R11903), .clock(clock), .in1(R11902));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11945 (.out1(R11946), .clock(clock), .in1(R11945));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12035 (.out1(R12036), .clock(clock), .in1(R12035));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12070 (.out1(R12071), .clock(clock), .in1(R12070));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12100 (.out1(R12101), .clock(clock), .in1(R12100));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12176 (.out1(R12177), .clock(clock), .in1(_1541));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12177 (.out1(R12178), .clock(clock), .in1(_1622));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1675 (.out1(_1623), .in1(R12178));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1676 (.out1(_1624), .in1(R12177), .in2(_1623));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1677 (.out1(idx_3674), .in1(_1624), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3911 (.out1(R3912), .clock(clock), .in1(R3911));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4167 (.out1(R4168), .clock(clock), .in1(R4167));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4422 (.out1(R4423), .clock(clock), .in1(R4422));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4667 (.out1(R4668), .clock(clock), .in1(R4667));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4907 (.out1(R4908), .clock(clock), .in1(R4907));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5194 (.out1(R5195), .clock(clock), .in1(R5194));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5426 (.out1(R5427), .clock(clock), .in1(R5426));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5653 (.out1(R5654), .clock(clock), .in1(R5653));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5927 (.out1(R5928), .clock(clock), .in1(R5927));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6145 (.out1(R6146), .clock(clock), .in1(R6145));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6358 (.out1(R6359), .clock(clock), .in1(R6358));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6619 (.out1(R6620), .clock(clock), .in1(R6619));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6824 (.out1(R6825), .clock(clock), .in1(R6824));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7024 (.out1(R7025), .clock(clock), .in1(R7024));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7271 (.out1(R7272), .clock(clock), .in1(R7271));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7463 (.out1(R7464), .clock(clock), .in1(R7463));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7650 (.out1(R7651), .clock(clock), .in1(R7650));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7884 (.out1(R7885), .clock(clock), .in1(R7884));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8063 (.out1(R8064), .clock(clock), .in1(R8063));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8237 (.out1(R8238), .clock(clock), .in1(R8237));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8458 (.out1(R8459), .clock(clock), .in1(R8458));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8624 (.out1(R8625), .clock(clock), .in1(R8624));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8785 (.out1(R8786), .clock(clock), .in1(R8785));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8993 (.out1(R8994), .clock(clock), .in1(R8993));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9146 (.out1(R9147), .clock(clock), .in1(R9146));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9294 (.out1(R9295), .clock(clock), .in1(R9294));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9489 (.out1(R9490), .clock(clock), .in1(R9489));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9629 (.out1(R9630), .clock(clock), .in1(R9629));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9764 (.out1(R9765), .clock(clock), .in1(R9764));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9946 (.out1(R9947), .clock(clock), .in1(R9946));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10073 (.out1(R10074), .clock(clock), .in1(R10073));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10195 (.out1(R10196), .clock(clock), .in1(R10195));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10364 (.out1(R10365), .clock(clock), .in1(R10364));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10477 (.out1(R10478), .clock(clock), .in1(R10477));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10585 (.out1(R10586), .clock(clock), .in1(R10585));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10741 (.out1(R10742), .clock(clock), .in1(R10741));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10841 (.out1(R10842), .clock(clock), .in1(R10841));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10936 (.out1(R10937), .clock(clock), .in1(R10936));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11078 (.out1(R11079), .clock(clock), .in1(R11078));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11165 (.out1(R11166), .clock(clock), .in1(R11165));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11247 (.out1(R11248), .clock(clock), .in1(R11247));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11376 (.out1(R11377), .clock(clock), .in1(R11376));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11450 (.out1(R11451), .clock(clock), .in1(R11450));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11519 (.out1(R11520), .clock(clock), .in1(R11519));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11635 (.out1(R11636), .clock(clock), .in1(R11635));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11696 (.out1(R11697), .clock(clock), .in1(R11696));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11752 (.out1(R11753), .clock(clock), .in1(R11752));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11855 (.out1(R11856), .clock(clock), .in1(R11855));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11903 (.out1(R11904), .clock(clock), .in1(R11903));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11946 (.out1(R11947), .clock(clock), .in1(R11946));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12036 (.out1(R12037), .clock(clock), .in1(R12036));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12071 (.out1(R12072), .clock(clock), .in1(R12071));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12101 (.out1(R12102), .clock(clock), .in1(R12101));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12178 (.out1(R12179), .clock(clock), .in1(idx_3674));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1681 (.out1(_1627), .in1(R12179));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1682 (.out1(_1628), .in1(_1627), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3912 (.out1(R3913), .clock(clock), .in1(R3912));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4168 (.out1(R4169), .clock(clock), .in1(R4168));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4423 (.out1(R4424), .clock(clock), .in1(R4423));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4668 (.out1(R4669), .clock(clock), .in1(R4668));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4908 (.out1(R4909), .clock(clock), .in1(R4908));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5195 (.out1(R5196), .clock(clock), .in1(R5195));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5427 (.out1(R5428), .clock(clock), .in1(R5427));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5654 (.out1(R5655), .clock(clock), .in1(R5654));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5928 (.out1(R5929), .clock(clock), .in1(R5928));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6146 (.out1(R6147), .clock(clock), .in1(R6146));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6359 (.out1(R6360), .clock(clock), .in1(R6359));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6620 (.out1(R6621), .clock(clock), .in1(R6620));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6825 (.out1(R6826), .clock(clock), .in1(R6825));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7025 (.out1(R7026), .clock(clock), .in1(R7025));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7272 (.out1(R7273), .clock(clock), .in1(R7272));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7464 (.out1(R7465), .clock(clock), .in1(R7464));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7651 (.out1(R7652), .clock(clock), .in1(R7651));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7885 (.out1(R7886), .clock(clock), .in1(R7885));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8064 (.out1(R8065), .clock(clock), .in1(R8064));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8238 (.out1(R8239), .clock(clock), .in1(R8238));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8459 (.out1(R8460), .clock(clock), .in1(R8459));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8625 (.out1(R8626), .clock(clock), .in1(R8625));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8786 (.out1(R8787), .clock(clock), .in1(R8786));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8994 (.out1(R8995), .clock(clock), .in1(R8994));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9147 (.out1(R9148), .clock(clock), .in1(R9147));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9295 (.out1(R9296), .clock(clock), .in1(R9295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9490 (.out1(R9491), .clock(clock), .in1(R9490));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9630 (.out1(R9631), .clock(clock), .in1(R9630));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9765 (.out1(R9766), .clock(clock), .in1(R9765));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9947 (.out1(R9948), .clock(clock), .in1(R9947));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10074 (.out1(R10075), .clock(clock), .in1(R10074));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10196 (.out1(R10197), .clock(clock), .in1(R10196));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10365 (.out1(R10366), .clock(clock), .in1(R10365));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10478 (.out1(R10479), .clock(clock), .in1(R10478));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10586 (.out1(R10587), .clock(clock), .in1(R10586));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10742 (.out1(R10743), .clock(clock), .in1(R10742));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10842 (.out1(R10843), .clock(clock), .in1(R10842));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10937 (.out1(R10938), .clock(clock), .in1(R10937));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11079 (.out1(R11080), .clock(clock), .in1(R11079));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11166 (.out1(R11167), .clock(clock), .in1(R11166));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11248 (.out1(R11249), .clock(clock), .in1(R11248));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11377 (.out1(R11378), .clock(clock), .in1(R11377));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11451 (.out1(R11452), .clock(clock), .in1(R11451));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11520 (.out1(R11521), .clock(clock), .in1(R11520));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11636 (.out1(R11637), .clock(clock), .in1(R11636));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11697 (.out1(R11698), .clock(clock), .in1(R11697));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11753 (.out1(R11754), .clock(clock), .in1(R11753));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11856 (.out1(R11857), .clock(clock), .in1(R11856));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11904 (.out1(R11905), .clock(clock), .in1(R11904));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11947 (.out1(R11948), .clock(clock), .in1(R11947));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12037 (.out1(R12038), .clock(clock), .in1(R12037));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12072 (.out1(R12073), .clock(clock), .in1(R12072));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12102 (.out1(R12103), .clock(clock), .in1(R12102));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12179 (.out1(R12180), .clock(clock), .in1(R12179));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12201 (.out1(R12202), .clock(clock), .in1(_1628));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1683 (.out1(_1629), .in1(vec118_3676_D), .in2(R12202));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3913 (.out1(R3914), .clock(clock), .in1(R3913));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4169 (.out1(R4170), .clock(clock), .in1(R4169));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4424 (.out1(R4425), .clock(clock), .in1(R4424));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4669 (.out1(R4670), .clock(clock), .in1(R4669));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4909 (.out1(R4910), .clock(clock), .in1(R4909));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5196 (.out1(R5197), .clock(clock), .in1(R5196));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5428 (.out1(R5429), .clock(clock), .in1(R5428));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5655 (.out1(R5656), .clock(clock), .in1(R5655));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5929 (.out1(R5930), .clock(clock), .in1(R5929));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6147 (.out1(R6148), .clock(clock), .in1(R6147));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6360 (.out1(R6361), .clock(clock), .in1(R6360));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6621 (.out1(R6622), .clock(clock), .in1(R6621));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6826 (.out1(R6827), .clock(clock), .in1(R6826));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7026 (.out1(R7027), .clock(clock), .in1(R7026));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7273 (.out1(R7274), .clock(clock), .in1(R7273));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7465 (.out1(R7466), .clock(clock), .in1(R7465));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7652 (.out1(R7653), .clock(clock), .in1(R7652));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7886 (.out1(R7887), .clock(clock), .in1(R7886));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8065 (.out1(R8066), .clock(clock), .in1(R8065));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8239 (.out1(R8240), .clock(clock), .in1(R8239));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8460 (.out1(R8461), .clock(clock), .in1(R8460));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8626 (.out1(R8627), .clock(clock), .in1(R8626));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8787 (.out1(R8788), .clock(clock), .in1(R8787));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8995 (.out1(R8996), .clock(clock), .in1(R8995));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9148 (.out1(R9149), .clock(clock), .in1(R9148));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9296 (.out1(R9297), .clock(clock), .in1(R9296));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9491 (.out1(R9492), .clock(clock), .in1(R9491));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9631 (.out1(R9632), .clock(clock), .in1(R9631));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9766 (.out1(R9767), .clock(clock), .in1(R9766));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9948 (.out1(R9949), .clock(clock), .in1(R9948));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10075 (.out1(R10076), .clock(clock), .in1(R10075));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10197 (.out1(R10198), .clock(clock), .in1(R10197));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10366 (.out1(R10367), .clock(clock), .in1(R10366));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10479 (.out1(R10480), .clock(clock), .in1(R10479));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10587 (.out1(R10588), .clock(clock), .in1(R10587));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10743 (.out1(R10744), .clock(clock), .in1(R10743));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10843 (.out1(R10844), .clock(clock), .in1(R10843));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10938 (.out1(R10939), .clock(clock), .in1(R10938));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11080 (.out1(R11081), .clock(clock), .in1(R11080));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11167 (.out1(R11168), .clock(clock), .in1(R11167));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11249 (.out1(R11250), .clock(clock), .in1(R11249));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11378 (.out1(R11379), .clock(clock), .in1(R11378));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11452 (.out1(R11453), .clock(clock), .in1(R11452));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11521 (.out1(R11522), .clock(clock), .in1(R11521));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11637 (.out1(R11638), .clock(clock), .in1(R11637));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11698 (.out1(R11699), .clock(clock), .in1(R11698));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11754 (.out1(R11755), .clock(clock), .in1(R11754));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11857 (.out1(R11858), .clock(clock), .in1(R11857));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11905 (.out1(R11906), .clock(clock), .in1(R11905));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11948 (.out1(R11949), .clock(clock), .in1(R11948));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12038 (.out1(R12039), .clock(clock), .in1(R12038));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12073 (.out1(R12074), .clock(clock), .in1(R12073));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12103 (.out1(R12104), .clock(clock), .in1(R12103));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12180 (.out1(R12181), .clock(clock), .in1(R12180));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12202 (.out1(R12203), .clock(clock), .in1(_1629));
  SRAM op1684 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1630),.ADR(R12203));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3914 (.out1(R3915), .clock(clock), .in1(R3914));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4170 (.out1(R4171), .clock(clock), .in1(R4170));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4425 (.out1(R4426), .clock(clock), .in1(R4425));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4670 (.out1(R4671), .clock(clock), .in1(R4670));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4910 (.out1(R4911), .clock(clock), .in1(R4910));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5197 (.out1(R5198), .clock(clock), .in1(R5197));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5429 (.out1(R5430), .clock(clock), .in1(R5429));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5656 (.out1(R5657), .clock(clock), .in1(R5656));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5930 (.out1(R5931), .clock(clock), .in1(R5930));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6148 (.out1(R6149), .clock(clock), .in1(R6148));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6361 (.out1(R6362), .clock(clock), .in1(R6361));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6622 (.out1(R6623), .clock(clock), .in1(R6622));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6827 (.out1(R6828), .clock(clock), .in1(R6827));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7027 (.out1(R7028), .clock(clock), .in1(R7027));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7274 (.out1(R7275), .clock(clock), .in1(R7274));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7466 (.out1(R7467), .clock(clock), .in1(R7466));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7653 (.out1(R7654), .clock(clock), .in1(R7653));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7887 (.out1(R7888), .clock(clock), .in1(R7887));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8066 (.out1(R8067), .clock(clock), .in1(R8066));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8240 (.out1(R8241), .clock(clock), .in1(R8240));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8461 (.out1(R8462), .clock(clock), .in1(R8461));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8627 (.out1(R8628), .clock(clock), .in1(R8627));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8788 (.out1(R8789), .clock(clock), .in1(R8788));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8996 (.out1(R8997), .clock(clock), .in1(R8996));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9149 (.out1(R9150), .clock(clock), .in1(R9149));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9297 (.out1(R9298), .clock(clock), .in1(R9297));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9492 (.out1(R9493), .clock(clock), .in1(R9492));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9632 (.out1(R9633), .clock(clock), .in1(R9632));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9767 (.out1(R9768), .clock(clock), .in1(R9767));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9949 (.out1(R9950), .clock(clock), .in1(R9949));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10076 (.out1(R10077), .clock(clock), .in1(R10076));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10198 (.out1(R10199), .clock(clock), .in1(R10198));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10367 (.out1(R10368), .clock(clock), .in1(R10367));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10480 (.out1(R10481), .clock(clock), .in1(R10480));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10588 (.out1(R10589), .clock(clock), .in1(R10588));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10744 (.out1(R10745), .clock(clock), .in1(R10744));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10844 (.out1(R10845), .clock(clock), .in1(R10844));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10939 (.out1(R10940), .clock(clock), .in1(R10939));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11081 (.out1(R11082), .clock(clock), .in1(R11081));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11168 (.out1(R11169), .clock(clock), .in1(R11168));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11250 (.out1(R11251), .clock(clock), .in1(R11250));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11379 (.out1(R11380), .clock(clock), .in1(R11379));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11453 (.out1(R11454), .clock(clock), .in1(R11453));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11522 (.out1(R11523), .clock(clock), .in1(R11522));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11638 (.out1(R11639), .clock(clock), .in1(R11638));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11699 (.out1(R11700), .clock(clock), .in1(R11699));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11755 (.out1(R11756), .clock(clock), .in1(R11755));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11858 (.out1(R11859), .clock(clock), .in1(R11858));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11906 (.out1(R11907), .clock(clock), .in1(R11906));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11949 (.out1(R11950), .clock(clock), .in1(R11949));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12039 (.out1(R12040), .clock(clock), .in1(R12039));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12074 (.out1(R12075), .clock(clock), .in1(R12074));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12104 (.out1(R12105), .clock(clock), .in1(R12104));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12181 (.out1(R12182), .clock(clock), .in1(R12181));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12203 (.out1(R12204), .clock(clock), .in1(_1630));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op1678 (.out1(_1625), .in1(ip2_3602_D), .in2(3 'd 4));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1679 (.out1(_1626), .in1(_1625));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op1680 (.out1(off_3675), .in1(_1626), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1685 (.out1(_1631), .in1(R12204), .in2(off_3675));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3915 (.out1(R3916), .clock(clock), .in1(R3915));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4171 (.out1(R4172), .clock(clock), .in1(R4171));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4426 (.out1(R4427), .clock(clock), .in1(R4426));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4671 (.out1(R4672), .clock(clock), .in1(R4671));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4911 (.out1(R4912), .clock(clock), .in1(R4911));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5198 (.out1(R5199), .clock(clock), .in1(R5198));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5430 (.out1(R5431), .clock(clock), .in1(R5430));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5657 (.out1(R5658), .clock(clock), .in1(R5657));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5931 (.out1(R5932), .clock(clock), .in1(R5931));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6149 (.out1(R6150), .clock(clock), .in1(R6149));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6362 (.out1(R6363), .clock(clock), .in1(R6362));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6623 (.out1(R6624), .clock(clock), .in1(R6623));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6828 (.out1(R6829), .clock(clock), .in1(R6828));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7028 (.out1(R7029), .clock(clock), .in1(R7028));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7275 (.out1(R7276), .clock(clock), .in1(R7275));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7467 (.out1(R7468), .clock(clock), .in1(R7467));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7654 (.out1(R7655), .clock(clock), .in1(R7654));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7888 (.out1(R7889), .clock(clock), .in1(R7888));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8067 (.out1(R8068), .clock(clock), .in1(R8067));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8241 (.out1(R8242), .clock(clock), .in1(R8241));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8462 (.out1(R8463), .clock(clock), .in1(R8462));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8628 (.out1(R8629), .clock(clock), .in1(R8628));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8789 (.out1(R8790), .clock(clock), .in1(R8789));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8997 (.out1(R8998), .clock(clock), .in1(R8997));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9150 (.out1(R9151), .clock(clock), .in1(R9150));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9298 (.out1(R9299), .clock(clock), .in1(R9298));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9493 (.out1(R9494), .clock(clock), .in1(R9493));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9633 (.out1(R9634), .clock(clock), .in1(R9633));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9768 (.out1(R9769), .clock(clock), .in1(R9768));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9950 (.out1(R9951), .clock(clock), .in1(R9950));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10077 (.out1(R10078), .clock(clock), .in1(R10077));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10199 (.out1(R10200), .clock(clock), .in1(R10199));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10368 (.out1(R10369), .clock(clock), .in1(R10368));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10481 (.out1(R10482), .clock(clock), .in1(R10481));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10589 (.out1(R10590), .clock(clock), .in1(R10589));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10745 (.out1(R10746), .clock(clock), .in1(R10745));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10845 (.out1(R10846), .clock(clock), .in1(R10845));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10940 (.out1(R10941), .clock(clock), .in1(R10940));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11082 (.out1(R11083), .clock(clock), .in1(R11082));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11169 (.out1(R11170), .clock(clock), .in1(R11169));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11251 (.out1(R11252), .clock(clock), .in1(R11251));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11380 (.out1(R11381), .clock(clock), .in1(R11380));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11454 (.out1(R11455), .clock(clock), .in1(R11454));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11523 (.out1(R11524), .clock(clock), .in1(R11523));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11639 (.out1(R11640), .clock(clock), .in1(R11639));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11700 (.out1(R11701), .clock(clock), .in1(R11700));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11756 (.out1(R11757), .clock(clock), .in1(R11756));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11859 (.out1(R11860), .clock(clock), .in1(R11859));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11907 (.out1(R11908), .clock(clock), .in1(R11907));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11950 (.out1(R11951), .clock(clock), .in1(R11950));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12040 (.out1(R12041), .clock(clock), .in1(R12040));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12075 (.out1(R12076), .clock(clock), .in1(R12075));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12105 (.out1(R12106), .clock(clock), .in1(R12105));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12182 (.out1(R12183), .clock(clock), .in1(R12182));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12204 (.out1(R12205), .clock(clock), .in1(off_3675));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12221 (.out1(R12222), .clock(clock), .in1(_1631));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op1686 (.out1(_1632), .in1(R12222), .in2(1 'd 1));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op1687 (.out1(ifout1687), .in1(_1632), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1755 (.out1(_1700), .in1(R12183));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1748 (.out1(_1693), .in1(R12183));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1737 (.out1(_1682), .in1(R12183));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1717 (.out1(_1662), .in1(R12183));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1756 (.out1(_1701), .in1(_1700), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1749 (.out1(_1694), .in1(_1693), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1738 (.out1(_1683), .in1(_1682), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1718 (.out1(_1663), .in1(_1662), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3916 (.out1(R3917), .clock(clock), .in1(R3916));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4172 (.out1(R4173), .clock(clock), .in1(R4172));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4427 (.out1(R4428), .clock(clock), .in1(R4427));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4672 (.out1(R4673), .clock(clock), .in1(R4672));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4912 (.out1(R4913), .clock(clock), .in1(R4912));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5199 (.out1(R5200), .clock(clock), .in1(R5199));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5431 (.out1(R5432), .clock(clock), .in1(R5431));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5658 (.out1(R5659), .clock(clock), .in1(R5658));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5932 (.out1(R5933), .clock(clock), .in1(R5932));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6150 (.out1(R6151), .clock(clock), .in1(R6150));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6363 (.out1(R6364), .clock(clock), .in1(R6363));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6624 (.out1(R6625), .clock(clock), .in1(R6624));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6829 (.out1(R6830), .clock(clock), .in1(R6829));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7029 (.out1(R7030), .clock(clock), .in1(R7029));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7276 (.out1(R7277), .clock(clock), .in1(R7276));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7468 (.out1(R7469), .clock(clock), .in1(R7468));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7655 (.out1(R7656), .clock(clock), .in1(R7655));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7889 (.out1(R7890), .clock(clock), .in1(R7889));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8068 (.out1(R8069), .clock(clock), .in1(R8068));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8242 (.out1(R8243), .clock(clock), .in1(R8242));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8463 (.out1(R8464), .clock(clock), .in1(R8463));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8629 (.out1(R8630), .clock(clock), .in1(R8629));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8790 (.out1(R8791), .clock(clock), .in1(R8790));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8998 (.out1(R8999), .clock(clock), .in1(R8998));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9151 (.out1(R9152), .clock(clock), .in1(R9151));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9299 (.out1(R9300), .clock(clock), .in1(R9299));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9494 (.out1(R9495), .clock(clock), .in1(R9494));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9634 (.out1(R9635), .clock(clock), .in1(R9634));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9769 (.out1(R9770), .clock(clock), .in1(R9769));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9951 (.out1(R9952), .clock(clock), .in1(R9951));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10078 (.out1(R10079), .clock(clock), .in1(R10078));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10200 (.out1(R10201), .clock(clock), .in1(R10200));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10369 (.out1(R10370), .clock(clock), .in1(R10369));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10482 (.out1(R10483), .clock(clock), .in1(R10482));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10590 (.out1(R10591), .clock(clock), .in1(R10590));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10746 (.out1(R10747), .clock(clock), .in1(R10746));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10846 (.out1(R10847), .clock(clock), .in1(R10846));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10941 (.out1(R10942), .clock(clock), .in1(R10941));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11083 (.out1(R11084), .clock(clock), .in1(R11083));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11170 (.out1(R11171), .clock(clock), .in1(R11170));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11252 (.out1(R11253), .clock(clock), .in1(R11252));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11381 (.out1(R11382), .clock(clock), .in1(R11381));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11455 (.out1(R11456), .clock(clock), .in1(R11455));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11524 (.out1(R11525), .clock(clock), .in1(R11524));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11640 (.out1(R11641), .clock(clock), .in1(R11640));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11701 (.out1(R11702), .clock(clock), .in1(R11701));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11757 (.out1(R11758), .clock(clock), .in1(R11757));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11860 (.out1(R11861), .clock(clock), .in1(R11860));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11908 (.out1(R11909), .clock(clock), .in1(R11908));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11951 (.out1(R11952), .clock(clock), .in1(R11951));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12041 (.out1(R12042), .clock(clock), .in1(R12041));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12076 (.out1(R12077), .clock(clock), .in1(R12076));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12106 (.out1(R12107), .clock(clock), .in1(R12106));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12183 (.out1(R12184), .clock(clock), .in1(R12183));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12205 (.out1(R12206), .clock(clock), .in1(R12205));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12222 (.out1(R12223), .clock(clock), .in1(ifout1687));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12246 (.out1(R12247), .clock(clock), .in1(_1701));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12247 (.out1(R12248), .clock(clock), .in1(_1694));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12248 (.out1(R12249), .clock(clock), .in1(_1683));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12249 (.out1(R12250), .clock(clock), .in1(_1663));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1730 (.out1(_1675), .in1(R12184));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1710 (.out1(_1655), .in1(R12184));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1699 (.out1(_1644), .in1(R12184));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1692 (.out1(_1637), .in1(R12184));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1759 (.out1(_1704), .in1(2 'd 2), .in2(R12206));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1731 (.out1(_1676), .in1(_1675), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1711 (.out1(_1656), .in1(_1655), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1700 (.out1(_1645), .in1(_1644), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1693 (.out1(_1638), .in1(_1637), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1757 (.out1(_1702), .in1(vec118_3676_D), .in2(R12247));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1750 (.out1(_1695), .in1(vec118_3676_D), .in2(R12248));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1739 (.out1(_1684), .in1(vec118_3676_D), .in2(R12249));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1719 (.out1(_1664), .in1(vec118_3676_D), .in2(R12250));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3917 (.out1(R3918), .clock(clock), .in1(R3917));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4173 (.out1(R4174), .clock(clock), .in1(R4173));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4428 (.out1(R4429), .clock(clock), .in1(R4428));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4673 (.out1(R4674), .clock(clock), .in1(R4673));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4913 (.out1(R4914), .clock(clock), .in1(R4913));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5200 (.out1(R5201), .clock(clock), .in1(R5200));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5432 (.out1(R5433), .clock(clock), .in1(R5432));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5659 (.out1(R5660), .clock(clock), .in1(R5659));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5933 (.out1(R5934), .clock(clock), .in1(R5933));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6151 (.out1(R6152), .clock(clock), .in1(R6151));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6364 (.out1(R6365), .clock(clock), .in1(R6364));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6625 (.out1(R6626), .clock(clock), .in1(R6625));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6830 (.out1(R6831), .clock(clock), .in1(R6830));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7030 (.out1(R7031), .clock(clock), .in1(R7030));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7277 (.out1(R7278), .clock(clock), .in1(R7277));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7469 (.out1(R7470), .clock(clock), .in1(R7469));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7656 (.out1(R7657), .clock(clock), .in1(R7656));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7890 (.out1(R7891), .clock(clock), .in1(R7890));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8069 (.out1(R8070), .clock(clock), .in1(R8069));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8243 (.out1(R8244), .clock(clock), .in1(R8243));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8464 (.out1(R8465), .clock(clock), .in1(R8464));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8630 (.out1(R8631), .clock(clock), .in1(R8630));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8791 (.out1(R8792), .clock(clock), .in1(R8791));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8999 (.out1(R9000), .clock(clock), .in1(R8999));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9152 (.out1(R9153), .clock(clock), .in1(R9152));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9300 (.out1(R9301), .clock(clock), .in1(R9300));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9495 (.out1(R9496), .clock(clock), .in1(R9495));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9635 (.out1(R9636), .clock(clock), .in1(R9635));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9770 (.out1(R9771), .clock(clock), .in1(R9770));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9952 (.out1(R9953), .clock(clock), .in1(R9952));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10079 (.out1(R10080), .clock(clock), .in1(R10079));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10201 (.out1(R10202), .clock(clock), .in1(R10201));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10370 (.out1(R10371), .clock(clock), .in1(R10370));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10483 (.out1(R10484), .clock(clock), .in1(R10483));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10591 (.out1(R10592), .clock(clock), .in1(R10591));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10747 (.out1(R10748), .clock(clock), .in1(R10747));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10847 (.out1(R10848), .clock(clock), .in1(R10847));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10942 (.out1(R10943), .clock(clock), .in1(R10942));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11084 (.out1(R11085), .clock(clock), .in1(R11084));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11171 (.out1(R11172), .clock(clock), .in1(R11171));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11253 (.out1(R11254), .clock(clock), .in1(R11253));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11382 (.out1(R11383), .clock(clock), .in1(R11382));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11456 (.out1(R11457), .clock(clock), .in1(R11456));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11525 (.out1(R11526), .clock(clock), .in1(R11525));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11641 (.out1(R11642), .clock(clock), .in1(R11641));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11702 (.out1(R11703), .clock(clock), .in1(R11702));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11758 (.out1(R11759), .clock(clock), .in1(R11758));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11861 (.out1(R11862), .clock(clock), .in1(R11861));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11909 (.out1(R11910), .clock(clock), .in1(R11909));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11952 (.out1(R11953), .clock(clock), .in1(R11952));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12042 (.out1(R12043), .clock(clock), .in1(R12042));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12077 (.out1(R12078), .clock(clock), .in1(R12077));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12107 (.out1(R12108), .clock(clock), .in1(R12107));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12184 (.out1(R12185), .clock(clock), .in1(R12184));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12206 (.out1(R12207), .clock(clock), .in1(R12206));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12223 (.out1(R12224), .clock(clock), .in1(R12223));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12250 (.out1(R12251), .clock(clock), .in1(_1704));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12251 (.out1(R12252), .clock(clock), .in1(_1676));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12252 (.out1(R12253), .clock(clock), .in1(_1656));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12253 (.out1(R12254), .clock(clock), .in1(_1645));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12254 (.out1(R12255), .clock(clock), .in1(_1638));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12255 (.out1(R12256), .clock(clock), .in1(_1702));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12256 (.out1(R12257), .clock(clock), .in1(_1695));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12257 (.out1(R12258), .clock(clock), .in1(_1684));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12258 (.out1(R12259), .clock(clock), .in1(_1664));
  SRAM op1758 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1703),.ADR(R12256));
  SRAM op1751 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1696),.ADR(R12257));
  SRAM op1740 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1685),.ADR(R12258));
  SRAM op1720 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1665),.ADR(R12259));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1752 (.out1(_1697), .in1(2 'd 2), .in2(R12207));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1741 (.out1(_1686), .in1(2 'd 2), .in2(R12207));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1734 (.out1(_1679), .in1(2 'd 2), .in2(R12207));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1721 (.out1(_1666), .in1(2 'd 2), .in2(R12207));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1714 (.out1(_1659), .in1(2 'd 2), .in2(R12207));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1703 (.out1(_1648), .in1(2 'd 2), .in2(R12207));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1732 (.out1(_1677), .in1(vec118_3676_D), .in2(R12252));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1712 (.out1(_1657), .in1(vec118_3676_D), .in2(R12253));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1701 (.out1(_1646), .in1(vec118_3676_D), .in2(R12254));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1694 (.out1(_1639), .in1(vec118_3676_D), .in2(R12255));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1760 (.out1(_1705), .in1(R12251), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3918 (.out1(R3919), .clock(clock), .in1(R3918));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4174 (.out1(R4175), .clock(clock), .in1(R4174));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4429 (.out1(R4430), .clock(clock), .in1(R4429));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4674 (.out1(R4675), .clock(clock), .in1(R4674));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4914 (.out1(R4915), .clock(clock), .in1(R4914));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5201 (.out1(R5202), .clock(clock), .in1(R5201));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5433 (.out1(R5434), .clock(clock), .in1(R5433));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5660 (.out1(R5661), .clock(clock), .in1(R5660));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5934 (.out1(R5935), .clock(clock), .in1(R5934));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6152 (.out1(R6153), .clock(clock), .in1(R6152));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6365 (.out1(R6366), .clock(clock), .in1(R6365));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6626 (.out1(R6627), .clock(clock), .in1(R6626));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6831 (.out1(R6832), .clock(clock), .in1(R6831));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7031 (.out1(R7032), .clock(clock), .in1(R7031));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7278 (.out1(R7279), .clock(clock), .in1(R7278));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7470 (.out1(R7471), .clock(clock), .in1(R7470));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7657 (.out1(R7658), .clock(clock), .in1(R7657));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7891 (.out1(R7892), .clock(clock), .in1(R7891));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8070 (.out1(R8071), .clock(clock), .in1(R8070));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8244 (.out1(R8245), .clock(clock), .in1(R8244));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8465 (.out1(R8466), .clock(clock), .in1(R8465));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8631 (.out1(R8632), .clock(clock), .in1(R8631));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8792 (.out1(R8793), .clock(clock), .in1(R8792));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9000 (.out1(R9001), .clock(clock), .in1(R9000));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9153 (.out1(R9154), .clock(clock), .in1(R9153));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9301 (.out1(R9302), .clock(clock), .in1(R9301));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9496 (.out1(R9497), .clock(clock), .in1(R9496));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9636 (.out1(R9637), .clock(clock), .in1(R9636));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9771 (.out1(R9772), .clock(clock), .in1(R9771));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9953 (.out1(R9954), .clock(clock), .in1(R9953));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10080 (.out1(R10081), .clock(clock), .in1(R10080));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10202 (.out1(R10203), .clock(clock), .in1(R10202));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10371 (.out1(R10372), .clock(clock), .in1(R10371));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10484 (.out1(R10485), .clock(clock), .in1(R10484));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10592 (.out1(R10593), .clock(clock), .in1(R10592));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10748 (.out1(R10749), .clock(clock), .in1(R10748));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10848 (.out1(R10849), .clock(clock), .in1(R10848));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10943 (.out1(R10944), .clock(clock), .in1(R10943));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11085 (.out1(R11086), .clock(clock), .in1(R11085));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11172 (.out1(R11173), .clock(clock), .in1(R11172));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11254 (.out1(R11255), .clock(clock), .in1(R11254));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11383 (.out1(R11384), .clock(clock), .in1(R11383));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11457 (.out1(R11458), .clock(clock), .in1(R11457));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11526 (.out1(R11527), .clock(clock), .in1(R11526));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11642 (.out1(R11643), .clock(clock), .in1(R11642));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11703 (.out1(R11704), .clock(clock), .in1(R11703));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11759 (.out1(R11760), .clock(clock), .in1(R11759));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11862 (.out1(R11863), .clock(clock), .in1(R11862));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11910 (.out1(R11911), .clock(clock), .in1(R11910));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11953 (.out1(R11954), .clock(clock), .in1(R11953));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12043 (.out1(R12044), .clock(clock), .in1(R12043));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12078 (.out1(R12079), .clock(clock), .in1(R12078));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12108 (.out1(R12109), .clock(clock), .in1(R12108));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12185 (.out1(R12186), .clock(clock), .in1(R12185));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12207 (.out1(R12208), .clock(clock), .in1(R12207));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12224 (.out1(R12225), .clock(clock), .in1(R12224));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12259 (.out1(R12260), .clock(clock), .in1(_1703));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12260 (.out1(R12261), .clock(clock), .in1(_1696));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12261 (.out1(R12262), .clock(clock), .in1(_1685));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12262 (.out1(R12263), .clock(clock), .in1(_1665));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12263 (.out1(R12264), .clock(clock), .in1(_1697));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12264 (.out1(R12265), .clock(clock), .in1(_1686));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12265 (.out1(R12266), .clock(clock), .in1(_1679));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12266 (.out1(R12267), .clock(clock), .in1(_1666));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12267 (.out1(R12268), .clock(clock), .in1(_1659));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12268 (.out1(R12269), .clock(clock), .in1(_1648));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12269 (.out1(R12270), .clock(clock), .in1(_1677));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12270 (.out1(R12271), .clock(clock), .in1(_1657));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12271 (.out1(R12272), .clock(clock), .in1(_1646));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12272 (.out1(R12273), .clock(clock), .in1(_1639));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12273 (.out1(R12274), .clock(clock), .in1(_1705));
  SRAM op1733 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1678),.ADR(R12270));
  SRAM op1713 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1658),.ADR(R12271));
  SRAM op1702 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1647),.ADR(R12272));
  SRAM op1695 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1640),.ADR(R12273));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1761 (.out1(_1706), .in1(R12260), .in2(R12274));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1762 (.out1(_1707), .in1(_1706), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1753 (.out1(_1698), .in1(R12264), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1742 (.out1(_1687), .in1(R12265), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1722 (.out1(_1667), .in1(R12267), .in2(64 'd 18446744073709551615));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1696 (.out1(_1641), .in1(2 'd 2), .in2(R12208));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1763 (.out1(_1708), .in1(_1707), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1754 (.out1(_1699), .in1(R12261), .in2(_1698));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1743 (.out1(_1688), .in1(R12262), .in2(_1687));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1723 (.out1(_1668), .in1(R12263), .in2(_1667));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1764 (.out1(_1709), .in1(_1699), .in2(_1708));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1744 (.out1(_1689), .in1(_1688), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1735 (.out1(_1680), .in1(R12266), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1724 (.out1(_1669), .in1(_1668), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1715 (.out1(_1660), .in1(R12268), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1704 (.out1(_1649), .in1(R12269), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3919 (.out1(R3920), .clock(clock), .in1(R3919));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4175 (.out1(R4176), .clock(clock), .in1(R4175));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4430 (.out1(R4431), .clock(clock), .in1(R4430));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4675 (.out1(R4676), .clock(clock), .in1(R4675));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4915 (.out1(R4916), .clock(clock), .in1(R4915));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5202 (.out1(R5203), .clock(clock), .in1(R5202));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5434 (.out1(R5435), .clock(clock), .in1(R5434));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5661 (.out1(R5662), .clock(clock), .in1(R5661));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5935 (.out1(R5936), .clock(clock), .in1(R5935));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6153 (.out1(R6154), .clock(clock), .in1(R6153));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6366 (.out1(R6367), .clock(clock), .in1(R6366));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6627 (.out1(R6628), .clock(clock), .in1(R6627));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6832 (.out1(R6833), .clock(clock), .in1(R6832));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7032 (.out1(R7033), .clock(clock), .in1(R7032));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7279 (.out1(R7280), .clock(clock), .in1(R7279));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7471 (.out1(R7472), .clock(clock), .in1(R7471));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7658 (.out1(R7659), .clock(clock), .in1(R7658));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7892 (.out1(R7893), .clock(clock), .in1(R7892));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8071 (.out1(R8072), .clock(clock), .in1(R8071));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8245 (.out1(R8246), .clock(clock), .in1(R8245));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8466 (.out1(R8467), .clock(clock), .in1(R8466));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8632 (.out1(R8633), .clock(clock), .in1(R8632));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8793 (.out1(R8794), .clock(clock), .in1(R8793));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9001 (.out1(R9002), .clock(clock), .in1(R9001));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9154 (.out1(R9155), .clock(clock), .in1(R9154));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9302 (.out1(R9303), .clock(clock), .in1(R9302));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9497 (.out1(R9498), .clock(clock), .in1(R9497));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9637 (.out1(R9638), .clock(clock), .in1(R9637));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9772 (.out1(R9773), .clock(clock), .in1(R9772));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9954 (.out1(R9955), .clock(clock), .in1(R9954));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10081 (.out1(R10082), .clock(clock), .in1(R10081));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10203 (.out1(R10204), .clock(clock), .in1(R10203));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10372 (.out1(R10373), .clock(clock), .in1(R10372));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10485 (.out1(R10486), .clock(clock), .in1(R10485));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10593 (.out1(R10594), .clock(clock), .in1(R10593));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10749 (.out1(R10750), .clock(clock), .in1(R10749));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10849 (.out1(R10850), .clock(clock), .in1(R10849));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10944 (.out1(R10945), .clock(clock), .in1(R10944));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11086 (.out1(R11087), .clock(clock), .in1(R11086));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11173 (.out1(R11174), .clock(clock), .in1(R11173));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11255 (.out1(R11256), .clock(clock), .in1(R11255));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11384 (.out1(R11385), .clock(clock), .in1(R11384));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11458 (.out1(R11459), .clock(clock), .in1(R11458));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11527 (.out1(R11528), .clock(clock), .in1(R11527));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11643 (.out1(R11644), .clock(clock), .in1(R11643));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11704 (.out1(R11705), .clock(clock), .in1(R11704));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11760 (.out1(R11761), .clock(clock), .in1(R11760));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11863 (.out1(R11864), .clock(clock), .in1(R11863));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11911 (.out1(R11912), .clock(clock), .in1(R11911));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11954 (.out1(R11955), .clock(clock), .in1(R11954));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12044 (.out1(R12045), .clock(clock), .in1(R12044));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12079 (.out1(R12080), .clock(clock), .in1(R12079));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12109 (.out1(R12110), .clock(clock), .in1(R12109));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12186 (.out1(R12187), .clock(clock), .in1(R12186));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12208 (.out1(R12209), .clock(clock), .in1(R12208));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12225 (.out1(R12226), .clock(clock), .in1(R12225));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12274 (.out1(R12275), .clock(clock), .in1(_1678));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12275 (.out1(R12276), .clock(clock), .in1(_1658));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12276 (.out1(R12277), .clock(clock), .in1(_1647));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12277 (.out1(R12278), .clock(clock), .in1(_1640));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12278 (.out1(R12279), .clock(clock), .in1(_1641));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12279 (.out1(R12280), .clock(clock), .in1(_1709));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12280 (.out1(R12281), .clock(clock), .in1(_1689));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12281 (.out1(R12282), .clock(clock), .in1(_1680));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12282 (.out1(R12283), .clock(clock), .in1(_1669));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12283 (.out1(R12284), .clock(clock), .in1(_1660));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12284 (.out1(R12285), .clock(clock), .in1(_1649));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1745 (.out1(_1690), .in1(R12281), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1736 (.out1(_1681), .in1(R12275), .in2(R12282));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1705 (.out1(_1650), .in1(R12277), .in2(R12285));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1765 (.out1(_1710), .in1(R12280), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1746 (.out1(_1691), .in1(_1681), .in2(_1690));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1725 (.out1(_1670), .in1(R12283), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1716 (.out1(_1661), .in1(R12276), .in2(R12284));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1706 (.out1(_1651), .in1(_1650), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1697 (.out1(_1642), .in1(R12279), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1726 (.out1(_1671), .in1(_1661), .in2(_1670));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1766 (.out1(_1711), .in1(_1710), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1747 (.out1(_1692), .in1(_1691), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1707 (.out1(_1652), .in1(_1651), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1698 (.out1(_1643), .in1(R12278), .in2(_1642));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1767 (.out1(_1712), .in1(_1692), .in2(_1711));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1727 (.out1(_1672), .in1(_1671), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1708 (.out1(_1653), .in1(_1643), .in2(_1652));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3920 (.out1(R3921), .clock(clock), .in1(R3920));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4176 (.out1(R4177), .clock(clock), .in1(R4176));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4431 (.out1(R4432), .clock(clock), .in1(R4431));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4676 (.out1(R4677), .clock(clock), .in1(R4676));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4916 (.out1(R4917), .clock(clock), .in1(R4916));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5203 (.out1(R5204), .clock(clock), .in1(R5203));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5435 (.out1(R5436), .clock(clock), .in1(R5435));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5662 (.out1(R5663), .clock(clock), .in1(R5662));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5936 (.out1(R5937), .clock(clock), .in1(R5936));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6154 (.out1(R6155), .clock(clock), .in1(R6154));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6367 (.out1(R6368), .clock(clock), .in1(R6367));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6628 (.out1(R6629), .clock(clock), .in1(R6628));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6833 (.out1(R6834), .clock(clock), .in1(R6833));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7033 (.out1(R7034), .clock(clock), .in1(R7033));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7280 (.out1(R7281), .clock(clock), .in1(R7280));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7472 (.out1(R7473), .clock(clock), .in1(R7472));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7659 (.out1(R7660), .clock(clock), .in1(R7659));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7893 (.out1(R7894), .clock(clock), .in1(R7893));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8072 (.out1(R8073), .clock(clock), .in1(R8072));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8246 (.out1(R8247), .clock(clock), .in1(R8246));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8467 (.out1(R8468), .clock(clock), .in1(R8467));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8633 (.out1(R8634), .clock(clock), .in1(R8633));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8794 (.out1(R8795), .clock(clock), .in1(R8794));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9002 (.out1(R9003), .clock(clock), .in1(R9002));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9155 (.out1(R9156), .clock(clock), .in1(R9155));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9303 (.out1(R9304), .clock(clock), .in1(R9303));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9498 (.out1(R9499), .clock(clock), .in1(R9498));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9638 (.out1(R9639), .clock(clock), .in1(R9638));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9773 (.out1(R9774), .clock(clock), .in1(R9773));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9955 (.out1(R9956), .clock(clock), .in1(R9955));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10082 (.out1(R10083), .clock(clock), .in1(R10082));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10204 (.out1(R10205), .clock(clock), .in1(R10204));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10373 (.out1(R10374), .clock(clock), .in1(R10373));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10486 (.out1(R10487), .clock(clock), .in1(R10486));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10594 (.out1(R10595), .clock(clock), .in1(R10594));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10750 (.out1(R10751), .clock(clock), .in1(R10750));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10850 (.out1(R10851), .clock(clock), .in1(R10850));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10945 (.out1(R10946), .clock(clock), .in1(R10945));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11087 (.out1(R11088), .clock(clock), .in1(R11087));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11174 (.out1(R11175), .clock(clock), .in1(R11174));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11256 (.out1(R11257), .clock(clock), .in1(R11256));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11385 (.out1(R11386), .clock(clock), .in1(R11385));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11459 (.out1(R11460), .clock(clock), .in1(R11459));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11528 (.out1(R11529), .clock(clock), .in1(R11528));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11644 (.out1(R11645), .clock(clock), .in1(R11644));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11705 (.out1(R11706), .clock(clock), .in1(R11705));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11761 (.out1(R11762), .clock(clock), .in1(R11761));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11864 (.out1(R11865), .clock(clock), .in1(R11864));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11912 (.out1(R11913), .clock(clock), .in1(R11912));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11955 (.out1(R11956), .clock(clock), .in1(R11955));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12045 (.out1(R12046), .clock(clock), .in1(R12045));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12080 (.out1(R12081), .clock(clock), .in1(R12080));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12110 (.out1(R12111), .clock(clock), .in1(R12110));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12187 (.out1(R12188), .clock(clock), .in1(R12187));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12209 (.out1(R12210), .clock(clock), .in1(R12209));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12226 (.out1(R12227), .clock(clock), .in1(R12226));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12285 (.out1(R12286), .clock(clock), .in1(_1712));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12286 (.out1(R12287), .clock(clock), .in1(_1672));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12287 (.out1(R12288), .clock(clock), .in1(_1653));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1688 (.out1(_1633), .in1(R12188));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1728 (.out1(_1673), .in1(R12287), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1709 (.out1(_1654), .in1(R12288), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op1768 (.out1(_1713), .in1(R12286), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1729 (.out1(_1674), .in1(_1654), .in2(_1673));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1689 (.out1(_1634), .in1(_1633), .in2(2 'd 2));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1769 (.out1(_1714), .in1(_1674), .in2(_1713));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op1770 (.out1(_1715), .in1(_1714), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3921 (.out1(R3922), .clock(clock), .in1(R3921));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4177 (.out1(R4178), .clock(clock), .in1(R4177));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4432 (.out1(R4433), .clock(clock), .in1(R4432));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4677 (.out1(R4678), .clock(clock), .in1(R4677));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4917 (.out1(R4918), .clock(clock), .in1(R4917));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5204 (.out1(R5205), .clock(clock), .in1(R5204));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5436 (.out1(R5437), .clock(clock), .in1(R5436));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5663 (.out1(R5664), .clock(clock), .in1(R5663));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5937 (.out1(R5938), .clock(clock), .in1(R5937));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6155 (.out1(R6156), .clock(clock), .in1(R6155));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6368 (.out1(R6369), .clock(clock), .in1(R6368));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6629 (.out1(R6630), .clock(clock), .in1(R6629));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6834 (.out1(R6835), .clock(clock), .in1(R6834));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7034 (.out1(R7035), .clock(clock), .in1(R7034));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7281 (.out1(R7282), .clock(clock), .in1(R7281));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7473 (.out1(R7474), .clock(clock), .in1(R7473));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7660 (.out1(R7661), .clock(clock), .in1(R7660));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7894 (.out1(R7895), .clock(clock), .in1(R7894));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8073 (.out1(R8074), .clock(clock), .in1(R8073));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8247 (.out1(R8248), .clock(clock), .in1(R8247));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8468 (.out1(R8469), .clock(clock), .in1(R8468));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8634 (.out1(R8635), .clock(clock), .in1(R8634));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8795 (.out1(R8796), .clock(clock), .in1(R8795));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9003 (.out1(R9004), .clock(clock), .in1(R9003));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9156 (.out1(R9157), .clock(clock), .in1(R9156));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9304 (.out1(R9305), .clock(clock), .in1(R9304));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9499 (.out1(R9500), .clock(clock), .in1(R9499));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9639 (.out1(R9640), .clock(clock), .in1(R9639));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9774 (.out1(R9775), .clock(clock), .in1(R9774));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9956 (.out1(R9957), .clock(clock), .in1(R9956));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10083 (.out1(R10084), .clock(clock), .in1(R10083));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10205 (.out1(R10206), .clock(clock), .in1(R10205));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10374 (.out1(R10375), .clock(clock), .in1(R10374));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10487 (.out1(R10488), .clock(clock), .in1(R10487));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10595 (.out1(R10596), .clock(clock), .in1(R10595));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10751 (.out1(R10752), .clock(clock), .in1(R10751));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10851 (.out1(R10852), .clock(clock), .in1(R10851));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10946 (.out1(R10947), .clock(clock), .in1(R10946));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11088 (.out1(R11089), .clock(clock), .in1(R11088));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11175 (.out1(R11176), .clock(clock), .in1(R11175));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11257 (.out1(R11258), .clock(clock), .in1(R11257));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11386 (.out1(R11387), .clock(clock), .in1(R11386));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11460 (.out1(R11461), .clock(clock), .in1(R11460));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11529 (.out1(R11530), .clock(clock), .in1(R11529));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11645 (.out1(R11646), .clock(clock), .in1(R11645));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11706 (.out1(R11707), .clock(clock), .in1(R11706));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11762 (.out1(R11763), .clock(clock), .in1(R11762));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11865 (.out1(R11866), .clock(clock), .in1(R11865));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11913 (.out1(R11914), .clock(clock), .in1(R11913));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11956 (.out1(R11957), .clock(clock), .in1(R11956));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12046 (.out1(R12047), .clock(clock), .in1(R12046));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12081 (.out1(R12082), .clock(clock), .in1(R12081));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12111 (.out1(R12112), .clock(clock), .in1(R12111));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12188 (.out1(R12189), .clock(clock), .in1(R12188));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12210 (.out1(R12211), .clock(clock), .in1(R12210));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12227 (.out1(R12228), .clock(clock), .in1(R12227));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12288 (.out1(R12289), .clock(clock), .in1(_1634));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12289 (.out1(R12290), .clock(clock), .in1(_1715));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op1771 (.out1(_1716), .in1(R12290), .in2(57 'd 72340172838076673));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1690 (.out1(_1635), .in1(base0_118_3681_D), .in2(R12289));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3922 (.out1(R3923), .clock(clock), .in1(R3922));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4178 (.out1(R4179), .clock(clock), .in1(R4178));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4433 (.out1(R4434), .clock(clock), .in1(R4433));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4678 (.out1(R4679), .clock(clock), .in1(R4678));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4918 (.out1(R4919), .clock(clock), .in1(R4918));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5205 (.out1(R5206), .clock(clock), .in1(R5205));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5437 (.out1(R5438), .clock(clock), .in1(R5437));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5664 (.out1(R5665), .clock(clock), .in1(R5664));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5938 (.out1(R5939), .clock(clock), .in1(R5938));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6156 (.out1(R6157), .clock(clock), .in1(R6156));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6369 (.out1(R6370), .clock(clock), .in1(R6369));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6630 (.out1(R6631), .clock(clock), .in1(R6630));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6835 (.out1(R6836), .clock(clock), .in1(R6835));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7035 (.out1(R7036), .clock(clock), .in1(R7035));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7282 (.out1(R7283), .clock(clock), .in1(R7282));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7474 (.out1(R7475), .clock(clock), .in1(R7474));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7661 (.out1(R7662), .clock(clock), .in1(R7661));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7895 (.out1(R7896), .clock(clock), .in1(R7895));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8074 (.out1(R8075), .clock(clock), .in1(R8074));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8248 (.out1(R8249), .clock(clock), .in1(R8248));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8469 (.out1(R8470), .clock(clock), .in1(R8469));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8635 (.out1(R8636), .clock(clock), .in1(R8635));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8796 (.out1(R8797), .clock(clock), .in1(R8796));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9004 (.out1(R9005), .clock(clock), .in1(R9004));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9157 (.out1(R9158), .clock(clock), .in1(R9157));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9305 (.out1(R9306), .clock(clock), .in1(R9305));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9500 (.out1(R9501), .clock(clock), .in1(R9500));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9640 (.out1(R9641), .clock(clock), .in1(R9640));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9775 (.out1(R9776), .clock(clock), .in1(R9775));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9957 (.out1(R9958), .clock(clock), .in1(R9957));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10084 (.out1(R10085), .clock(clock), .in1(R10084));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10206 (.out1(R10207), .clock(clock), .in1(R10206));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10375 (.out1(R10376), .clock(clock), .in1(R10375));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10488 (.out1(R10489), .clock(clock), .in1(R10488));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10596 (.out1(R10597), .clock(clock), .in1(R10596));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10752 (.out1(R10753), .clock(clock), .in1(R10752));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10852 (.out1(R10853), .clock(clock), .in1(R10852));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10947 (.out1(R10948), .clock(clock), .in1(R10947));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11089 (.out1(R11090), .clock(clock), .in1(R11089));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11176 (.out1(R11177), .clock(clock), .in1(R11176));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11258 (.out1(R11259), .clock(clock), .in1(R11258));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11387 (.out1(R11388), .clock(clock), .in1(R11387));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11461 (.out1(R11462), .clock(clock), .in1(R11461));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11530 (.out1(R11531), .clock(clock), .in1(R11530));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11646 (.out1(R11647), .clock(clock), .in1(R11646));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11707 (.out1(R11708), .clock(clock), .in1(R11707));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11763 (.out1(R11764), .clock(clock), .in1(R11763));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11866 (.out1(R11867), .clock(clock), .in1(R11866));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11914 (.out1(R11915), .clock(clock), .in1(R11914));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11957 (.out1(R11958), .clock(clock), .in1(R11957));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12047 (.out1(R12048), .clock(clock), .in1(R12047));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12082 (.out1(R12083), .clock(clock), .in1(R12082));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12112 (.out1(R12113), .clock(clock), .in1(R12112));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12189 (.out1(R12190), .clock(clock), .in1(R12189));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12211 (.out1(R12212), .clock(clock), .in1(R12211));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12228 (.out1(R12229), .clock(clock), .in1(R12228));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12290 (.out1(R12291), .clock(clock), .in1(_1716));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12291 (.out1(R12292), .clock(clock), .in1(_1635));
  SRAM op1691 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1636),.ADR(R12292));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op1772 (.out1(_1717), .in1(R12291), .in2(6 'd 56));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3923 (.out1(R3924), .clock(clock), .in1(R3923));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4179 (.out1(R4180), .clock(clock), .in1(R4179));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4434 (.out1(R4435), .clock(clock), .in1(R4434));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4679 (.out1(R4680), .clock(clock), .in1(R4679));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4919 (.out1(R4920), .clock(clock), .in1(R4919));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5206 (.out1(R5207), .clock(clock), .in1(R5206));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5438 (.out1(R5439), .clock(clock), .in1(R5438));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5665 (.out1(R5666), .clock(clock), .in1(R5665));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5939 (.out1(R5940), .clock(clock), .in1(R5939));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6157 (.out1(R6158), .clock(clock), .in1(R6157));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6370 (.out1(R6371), .clock(clock), .in1(R6370));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6631 (.out1(R6632), .clock(clock), .in1(R6631));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6836 (.out1(R6837), .clock(clock), .in1(R6836));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7036 (.out1(R7037), .clock(clock), .in1(R7036));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7283 (.out1(R7284), .clock(clock), .in1(R7283));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7475 (.out1(R7476), .clock(clock), .in1(R7475));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7662 (.out1(R7663), .clock(clock), .in1(R7662));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7896 (.out1(R7897), .clock(clock), .in1(R7896));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8075 (.out1(R8076), .clock(clock), .in1(R8075));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8249 (.out1(R8250), .clock(clock), .in1(R8249));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8470 (.out1(R8471), .clock(clock), .in1(R8470));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8636 (.out1(R8637), .clock(clock), .in1(R8636));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8797 (.out1(R8798), .clock(clock), .in1(R8797));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9005 (.out1(R9006), .clock(clock), .in1(R9005));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9158 (.out1(R9159), .clock(clock), .in1(R9158));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9306 (.out1(R9307), .clock(clock), .in1(R9306));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9501 (.out1(R9502), .clock(clock), .in1(R9501));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9641 (.out1(R9642), .clock(clock), .in1(R9641));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9776 (.out1(R9777), .clock(clock), .in1(R9776));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9958 (.out1(R9959), .clock(clock), .in1(R9958));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10085 (.out1(R10086), .clock(clock), .in1(R10085));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10207 (.out1(R10208), .clock(clock), .in1(R10207));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10376 (.out1(R10377), .clock(clock), .in1(R10376));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10489 (.out1(R10490), .clock(clock), .in1(R10489));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10597 (.out1(R10598), .clock(clock), .in1(R10597));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10753 (.out1(R10754), .clock(clock), .in1(R10753));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10853 (.out1(R10854), .clock(clock), .in1(R10853));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10948 (.out1(R10949), .clock(clock), .in1(R10948));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11090 (.out1(R11091), .clock(clock), .in1(R11090));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11177 (.out1(R11178), .clock(clock), .in1(R11177));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11259 (.out1(R11260), .clock(clock), .in1(R11259));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11388 (.out1(R11389), .clock(clock), .in1(R11388));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11462 (.out1(R11463), .clock(clock), .in1(R11462));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11531 (.out1(R11532), .clock(clock), .in1(R11531));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11647 (.out1(R11648), .clock(clock), .in1(R11647));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11708 (.out1(R11709), .clock(clock), .in1(R11708));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11764 (.out1(R11765), .clock(clock), .in1(R11764));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11867 (.out1(R11868), .clock(clock), .in1(R11867));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11915 (.out1(R11916), .clock(clock), .in1(R11915));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11958 (.out1(R11959), .clock(clock), .in1(R11958));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12048 (.out1(R12049), .clock(clock), .in1(R12048));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12083 (.out1(R12084), .clock(clock), .in1(R12083));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12113 (.out1(R12114), .clock(clock), .in1(R12113));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12190 (.out1(R12191), .clock(clock), .in1(R12190));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12212 (.out1(R12213), .clock(clock), .in1(R12212));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12229 (.out1(R12230), .clock(clock), .in1(R12229));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12292 (.out1(R12293), .clock(clock), .in1(_1636));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12293 (.out1(R12294), .clock(clock), .in1(_1717));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1773 (.out1(_1718), .in1(R12294));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1774 (.out1(_1719), .in1(R12293), .in2(_1718));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1775 (.out1(idx_3682), .in1(_1719), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3924 (.out1(R3925), .clock(clock), .in1(R3924));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4180 (.out1(R4181), .clock(clock), .in1(R4180));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4435 (.out1(R4436), .clock(clock), .in1(R4435));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4680 (.out1(R4681), .clock(clock), .in1(R4680));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4920 (.out1(R4921), .clock(clock), .in1(R4920));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5207 (.out1(R5208), .clock(clock), .in1(R5207));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5439 (.out1(R5440), .clock(clock), .in1(R5439));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5666 (.out1(R5667), .clock(clock), .in1(R5666));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5940 (.out1(R5941), .clock(clock), .in1(R5940));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6158 (.out1(R6159), .clock(clock), .in1(R6158));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6371 (.out1(R6372), .clock(clock), .in1(R6371));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6632 (.out1(R6633), .clock(clock), .in1(R6632));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6837 (.out1(R6838), .clock(clock), .in1(R6837));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7037 (.out1(R7038), .clock(clock), .in1(R7037));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7284 (.out1(R7285), .clock(clock), .in1(R7284));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7476 (.out1(R7477), .clock(clock), .in1(R7476));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7663 (.out1(R7664), .clock(clock), .in1(R7663));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7897 (.out1(R7898), .clock(clock), .in1(R7897));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8076 (.out1(R8077), .clock(clock), .in1(R8076));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8250 (.out1(R8251), .clock(clock), .in1(R8250));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8471 (.out1(R8472), .clock(clock), .in1(R8471));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8637 (.out1(R8638), .clock(clock), .in1(R8637));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8798 (.out1(R8799), .clock(clock), .in1(R8798));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9006 (.out1(R9007), .clock(clock), .in1(R9006));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9159 (.out1(R9160), .clock(clock), .in1(R9159));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9307 (.out1(R9308), .clock(clock), .in1(R9307));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9502 (.out1(R9503), .clock(clock), .in1(R9502));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9642 (.out1(R9643), .clock(clock), .in1(R9642));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9777 (.out1(R9778), .clock(clock), .in1(R9777));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9959 (.out1(R9960), .clock(clock), .in1(R9959));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10086 (.out1(R10087), .clock(clock), .in1(R10086));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10208 (.out1(R10209), .clock(clock), .in1(R10208));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10377 (.out1(R10378), .clock(clock), .in1(R10377));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10490 (.out1(R10491), .clock(clock), .in1(R10490));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10598 (.out1(R10599), .clock(clock), .in1(R10598));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10754 (.out1(R10755), .clock(clock), .in1(R10754));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10854 (.out1(R10855), .clock(clock), .in1(R10854));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10949 (.out1(R10950), .clock(clock), .in1(R10949));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11091 (.out1(R11092), .clock(clock), .in1(R11091));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11178 (.out1(R11179), .clock(clock), .in1(R11178));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11260 (.out1(R11261), .clock(clock), .in1(R11260));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11389 (.out1(R11390), .clock(clock), .in1(R11389));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11463 (.out1(R11464), .clock(clock), .in1(R11463));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11532 (.out1(R11533), .clock(clock), .in1(R11532));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11648 (.out1(R11649), .clock(clock), .in1(R11648));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11709 (.out1(R11710), .clock(clock), .in1(R11709));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11765 (.out1(R11766), .clock(clock), .in1(R11765));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11868 (.out1(R11869), .clock(clock), .in1(R11868));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11916 (.out1(R11917), .clock(clock), .in1(R11916));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11959 (.out1(R11960), .clock(clock), .in1(R11959));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12049 (.out1(R12050), .clock(clock), .in1(R12049));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12084 (.out1(R12085), .clock(clock), .in1(R12084));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12114 (.out1(R12115), .clock(clock), .in1(R12114));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12191 (.out1(R12192), .clock(clock), .in1(R12191));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12213 (.out1(R12214), .clock(clock), .in1(R12213));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12230 (.out1(R12231), .clock(clock), .in1(R12230));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12294 (.out1(R12295), .clock(clock), .in1(idx_3682));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2563 (.out1(_2482), .in1(R10378));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2465 (.out1(_2387), .in1(R10755));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2367 (.out1(_2292), .in1(R11092));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2269 (.out1(_2197), .in1(R11390));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2171 (.out1(_2102), .in1(R11649));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2073 (.out1(_2007), .in1(R11869));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1975 (.out1(_1912), .in1(R12050));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1877 (.out1(_1817), .in1(R12192));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1779 (.out1(_1722), .in1(R12295));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2564 (.out1(_2483), .in1(_2482), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2466 (.out1(_2388), .in1(_2387), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2368 (.out1(_2293), .in1(_2292), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2270 (.out1(_2198), .in1(_2197), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2172 (.out1(_2103), .in1(_2102), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2074 (.out1(_2008), .in1(_2007), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1976 (.out1(_1913), .in1(_1912), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1878 (.out1(_1818), .in1(_1817), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1780 (.out1(_1723), .in1(_1722), .in2(2 'd 3));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3925 (.out1(R3926), .clock(clock), .in1(R3925));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4181 (.out1(R4182), .clock(clock), .in1(R4181));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4436 (.out1(R4437), .clock(clock), .in1(R4436));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4681 (.out1(R4682), .clock(clock), .in1(R4681));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4921 (.out1(R4922), .clock(clock), .in1(R4921));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5208 (.out1(R5209), .clock(clock), .in1(R5208));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5440 (.out1(R5441), .clock(clock), .in1(R5440));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5667 (.out1(R5668), .clock(clock), .in1(R5667));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5941 (.out1(R5942), .clock(clock), .in1(R5941));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6159 (.out1(R6160), .clock(clock), .in1(R6159));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6372 (.out1(R6373), .clock(clock), .in1(R6372));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6633 (.out1(R6634), .clock(clock), .in1(R6633));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6838 (.out1(R6839), .clock(clock), .in1(R6838));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7038 (.out1(R7039), .clock(clock), .in1(R7038));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7285 (.out1(R7286), .clock(clock), .in1(R7285));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7477 (.out1(R7478), .clock(clock), .in1(R7477));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7664 (.out1(R7665), .clock(clock), .in1(R7664));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7898 (.out1(R7899), .clock(clock), .in1(R7898));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8077 (.out1(R8078), .clock(clock), .in1(R8077));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8251 (.out1(R8252), .clock(clock), .in1(R8251));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8472 (.out1(R8473), .clock(clock), .in1(R8472));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8638 (.out1(R8639), .clock(clock), .in1(R8638));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8799 (.out1(R8800), .clock(clock), .in1(R8799));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9007 (.out1(R9008), .clock(clock), .in1(R9007));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9160 (.out1(R9161), .clock(clock), .in1(R9160));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9308 (.out1(R9309), .clock(clock), .in1(R9308));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9503 (.out1(R9504), .clock(clock), .in1(R9503));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9643 (.out1(R9644), .clock(clock), .in1(R9643));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9778 (.out1(R9779), .clock(clock), .in1(R9778));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9960 (.out1(R9961), .clock(clock), .in1(R9960));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10087 (.out1(R10088), .clock(clock), .in1(R10087));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10209 (.out1(R10210), .clock(clock), .in1(R10209));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10378 (.out1(R10379), .clock(clock), .in1(R10378));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10491 (.out1(R10492), .clock(clock), .in1(R10491));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10599 (.out1(R10600), .clock(clock), .in1(R10599));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10755 (.out1(R10756), .clock(clock), .in1(R10755));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10855 (.out1(R10856), .clock(clock), .in1(R10855));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10950 (.out1(R10951), .clock(clock), .in1(R10950));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11092 (.out1(R11093), .clock(clock), .in1(R11092));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11179 (.out1(R11180), .clock(clock), .in1(R11179));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11261 (.out1(R11262), .clock(clock), .in1(R11261));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11390 (.out1(R11391), .clock(clock), .in1(R11390));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11464 (.out1(R11465), .clock(clock), .in1(R11464));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11533 (.out1(R11534), .clock(clock), .in1(R11533));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11649 (.out1(R11650), .clock(clock), .in1(R11649));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11710 (.out1(R11711), .clock(clock), .in1(R11710));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11766 (.out1(R11767), .clock(clock), .in1(R11766));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11869 (.out1(R11870), .clock(clock), .in1(R11869));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11917 (.out1(R11918), .clock(clock), .in1(R11917));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11960 (.out1(R11961), .clock(clock), .in1(R11960));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12050 (.out1(R12051), .clock(clock), .in1(R12050));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12085 (.out1(R12086), .clock(clock), .in1(R12085));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12115 (.out1(R12116), .clock(clock), .in1(R12115));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12192 (.out1(R12193), .clock(clock), .in1(R12192));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12214 (.out1(R12215), .clock(clock), .in1(R12214));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12231 (.out1(R12232), .clock(clock), .in1(R12231));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12295 (.out1(R12296), .clock(clock), .in1(R12295));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12304 (.out1(R12305), .clock(clock), .in1(_2483));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12305 (.out1(R12306), .clock(clock), .in1(_2388));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12306 (.out1(R12307), .clock(clock), .in1(_2293));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12307 (.out1(R12308), .clock(clock), .in1(_2198));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12308 (.out1(R12309), .clock(clock), .in1(_2103));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12309 (.out1(R12310), .clock(clock), .in1(_2008));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12310 (.out1(R12311), .clock(clock), .in1(_1913));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12311 (.out1(R12312), .clock(clock), .in1(_1818));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12312 (.out1(R12313), .clock(clock), .in1(_1723));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3347 (.out1(_3242), .in1(R5942));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3249 (.out1(_3147), .in1(R6634));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3151 (.out1(_3052), .in1(R7286));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3053 (.out1(_2957), .in1(R7899));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2955 (.out1(_2862), .in1(R8473));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2857 (.out1(_2767), .in1(R9008));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2759 (.out1(_2672), .in1(R9504));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2661 (.out1(_2577), .in1(R9961));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3348 (.out1(_3243), .in1(_3242), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3250 (.out1(_3148), .in1(_3147), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3152 (.out1(_3053), .in1(_3052), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3054 (.out1(_2958), .in1(_2957), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2956 (.out1(_2863), .in1(_2862), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2858 (.out1(_2768), .in1(_2767), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2760 (.out1(_2673), .in1(_2672), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2662 (.out1(_2578), .in1(_2577), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2565 (.out1(_2484), .in1(leafvec76_3621_D), .in2(R12305));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2467 (.out1(_2389), .in1(leafvec82_3629_D), .in2(R12306));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2369 (.out1(_2294), .in1(leafvec88_3637_D), .in2(R12307));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2271 (.out1(_2199), .in1(leafvec94_3645_D), .in2(R12308));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2173 (.out1(_2104), .in1(leafvec100_3653_D), .in2(R12309));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2075 (.out1(_2009), .in1(leafvec106_3661_D), .in2(R12310));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1977 (.out1(_1914), .in1(leafvec112_3669_D), .in2(R12311));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1879 (.out1(_1819), .in1(leafvec118_3677_D), .in2(R12312));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1781 (.out1(_1724), .in1(leafvec124_3684_D), .in2(R12313));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3926 (.out1(R3927), .clock(clock), .in1(R3926));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4182 (.out1(R4183), .clock(clock), .in1(R4182));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4437 (.out1(R4438), .clock(clock), .in1(R4437));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4682 (.out1(R4683), .clock(clock), .in1(R4682));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4922 (.out1(R4923), .clock(clock), .in1(R4922));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5209 (.out1(R5210), .clock(clock), .in1(R5209));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5441 (.out1(R5442), .clock(clock), .in1(R5441));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5668 (.out1(R5669), .clock(clock), .in1(R5668));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5942 (.out1(R5943), .clock(clock), .in1(R5942));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6160 (.out1(R6161), .clock(clock), .in1(R6160));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6373 (.out1(R6374), .clock(clock), .in1(R6373));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6634 (.out1(R6635), .clock(clock), .in1(R6634));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6839 (.out1(R6840), .clock(clock), .in1(R6839));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7039 (.out1(R7040), .clock(clock), .in1(R7039));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7286 (.out1(R7287), .clock(clock), .in1(R7286));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7478 (.out1(R7479), .clock(clock), .in1(R7478));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7665 (.out1(R7666), .clock(clock), .in1(R7665));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7899 (.out1(R7900), .clock(clock), .in1(R7899));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8078 (.out1(R8079), .clock(clock), .in1(R8078));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8252 (.out1(R8253), .clock(clock), .in1(R8252));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8473 (.out1(R8474), .clock(clock), .in1(R8473));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8639 (.out1(R8640), .clock(clock), .in1(R8639));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8800 (.out1(R8801), .clock(clock), .in1(R8800));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9008 (.out1(R9009), .clock(clock), .in1(R9008));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9161 (.out1(R9162), .clock(clock), .in1(R9161));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9309 (.out1(R9310), .clock(clock), .in1(R9309));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9504 (.out1(R9505), .clock(clock), .in1(R9504));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9644 (.out1(R9645), .clock(clock), .in1(R9644));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9779 (.out1(R9780), .clock(clock), .in1(R9779));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9961 (.out1(R9962), .clock(clock), .in1(R9961));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10088 (.out1(R10089), .clock(clock), .in1(R10088));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10210 (.out1(R10211), .clock(clock), .in1(R10210));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10379 (.out1(R10380), .clock(clock), .in1(R10379));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10492 (.out1(R10493), .clock(clock), .in1(R10492));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10600 (.out1(R10601), .clock(clock), .in1(R10600));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10756 (.out1(R10757), .clock(clock), .in1(R10756));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10856 (.out1(R10857), .clock(clock), .in1(R10856));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10951 (.out1(R10952), .clock(clock), .in1(R10951));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11093 (.out1(R11094), .clock(clock), .in1(R11093));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11180 (.out1(R11181), .clock(clock), .in1(R11180));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11262 (.out1(R11263), .clock(clock), .in1(R11262));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11391 (.out1(R11392), .clock(clock), .in1(R11391));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11465 (.out1(R11466), .clock(clock), .in1(R11465));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11534 (.out1(R11535), .clock(clock), .in1(R11534));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11650 (.out1(R11651), .clock(clock), .in1(R11650));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11711 (.out1(R11712), .clock(clock), .in1(R11711));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11767 (.out1(R11768), .clock(clock), .in1(R11767));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11870 (.out1(R11871), .clock(clock), .in1(R11870));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11918 (.out1(R11919), .clock(clock), .in1(R11918));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11961 (.out1(R11962), .clock(clock), .in1(R11961));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12051 (.out1(R12052), .clock(clock), .in1(R12051));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12086 (.out1(R12087), .clock(clock), .in1(R12086));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12116 (.out1(R12117), .clock(clock), .in1(R12116));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12193 (.out1(R12194), .clock(clock), .in1(R12193));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12215 (.out1(R12216), .clock(clock), .in1(R12215));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12232 (.out1(R12233), .clock(clock), .in1(R12232));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12296 (.out1(R12297), .clock(clock), .in1(R12296));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12313 (.out1(R12314), .clock(clock), .in1(_3243));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12314 (.out1(R12315), .clock(clock), .in1(_3148));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12315 (.out1(R12316), .clock(clock), .in1(_3053));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12316 (.out1(R12317), .clock(clock), .in1(_2958));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12317 (.out1(R12318), .clock(clock), .in1(_2863));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12318 (.out1(R12319), .clock(clock), .in1(_2768));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12319 (.out1(R12320), .clock(clock), .in1(_2673));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12320 (.out1(R12321), .clock(clock), .in1(_2578));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12321 (.out1(R12322), .clock(clock), .in1(_2484));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12322 (.out1(R12323), .clock(clock), .in1(_2389));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12323 (.out1(R12324), .clock(clock), .in1(_2294));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12324 (.out1(R12325), .clock(clock), .in1(_2199));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12325 (.out1(R12326), .clock(clock), .in1(_2104));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12326 (.out1(R12327), .clock(clock), .in1(_2009));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12327 (.out1(R12328), .clock(clock), .in1(_1914));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12328 (.out1(R12329), .clock(clock), .in1(_1819));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12329 (.out1(R12330), .clock(clock), .in1(_1724));
  SRAM op2566 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2485),.ADR(R12322));
  SRAM op2468 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2390),.ADR(R12323));
  SRAM op2370 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2295),.ADR(R12324));
  SRAM op2272 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2200),.ADR(R12325));
  SRAM op2174 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2105),.ADR(R12326));
  SRAM op2076 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2010),.ADR(R12327));
  SRAM op1978 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1915),.ADR(R12328));
  SRAM op1880 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1820),.ADR(R12329));
  SRAM op1782 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1725),.ADR(R12330));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3543 (.out1(_3432), .in1(R4438));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3445 (.out1(_3337), .in1(R5210));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3544 (.out1(_3433), .in1(_3432), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3446 (.out1(_3338), .in1(_3337), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1776 (.out1(_1720), .in1(ip2_3602_D), .in2(2 'd 2));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3349 (.out1(_3244), .in1(leafvec28_3556_D), .in2(R12314));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3251 (.out1(_3149), .in1(leafvec34_3564_D), .in2(R12315));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3153 (.out1(_3054), .in1(leafvec40_3572_D), .in2(R12316));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3055 (.out1(_2959), .in1(leafvec46_3580_D), .in2(R12317));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2957 (.out1(_2864), .in1(leafvec52_3588_D), .in2(R12318));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2859 (.out1(_2769), .in1(leafvec58_3596_D), .in2(R12319));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2761 (.out1(_2674), .in1(leafvec64_3605_D), .in2(R12320));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2663 (.out1(_2579), .in1(leafvec70_3613_D), .in2(R12321));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3927 (.out1(R3928), .clock(clock), .in1(R3927));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4183 (.out1(R4184), .clock(clock), .in1(R4183));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4438 (.out1(R4439), .clock(clock), .in1(R4438));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4683 (.out1(R4684), .clock(clock), .in1(R4683));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4923 (.out1(R4924), .clock(clock), .in1(R4923));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5210 (.out1(R5211), .clock(clock), .in1(R5210));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5442 (.out1(R5443), .clock(clock), .in1(R5442));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5669 (.out1(R5670), .clock(clock), .in1(R5669));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5943 (.out1(R5944), .clock(clock), .in1(R5943));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6161 (.out1(R6162), .clock(clock), .in1(R6161));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6374 (.out1(R6375), .clock(clock), .in1(R6374));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6635 (.out1(R6636), .clock(clock), .in1(R6635));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6840 (.out1(R6841), .clock(clock), .in1(R6840));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7040 (.out1(R7041), .clock(clock), .in1(R7040));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7287 (.out1(R7288), .clock(clock), .in1(R7287));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7479 (.out1(R7480), .clock(clock), .in1(R7479));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7666 (.out1(R7667), .clock(clock), .in1(R7666));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7900 (.out1(R7901), .clock(clock), .in1(R7900));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8079 (.out1(R8080), .clock(clock), .in1(R8079));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8253 (.out1(R8254), .clock(clock), .in1(R8253));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8474 (.out1(R8475), .clock(clock), .in1(R8474));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8640 (.out1(R8641), .clock(clock), .in1(R8640));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8801 (.out1(R8802), .clock(clock), .in1(R8801));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9009 (.out1(R9010), .clock(clock), .in1(R9009));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9162 (.out1(R9163), .clock(clock), .in1(R9162));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9310 (.out1(R9311), .clock(clock), .in1(R9310));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9505 (.out1(R9506), .clock(clock), .in1(R9505));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9645 (.out1(R9646), .clock(clock), .in1(R9645));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9780 (.out1(R9781), .clock(clock), .in1(R9780));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9962 (.out1(R9963), .clock(clock), .in1(R9962));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10089 (.out1(R10090), .clock(clock), .in1(R10089));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10211 (.out1(R10212), .clock(clock), .in1(R10211));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10380 (.out1(R10381), .clock(clock), .in1(R10380));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10493 (.out1(R10494), .clock(clock), .in1(R10493));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10601 (.out1(R10602), .clock(clock), .in1(R10601));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10757 (.out1(R10758), .clock(clock), .in1(R10757));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10857 (.out1(R10858), .clock(clock), .in1(R10857));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10952 (.out1(R10953), .clock(clock), .in1(R10952));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11094 (.out1(R11095), .clock(clock), .in1(R11094));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11181 (.out1(R11182), .clock(clock), .in1(R11181));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11263 (.out1(R11264), .clock(clock), .in1(R11263));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11392 (.out1(R11393), .clock(clock), .in1(R11392));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11466 (.out1(R11467), .clock(clock), .in1(R11466));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11535 (.out1(R11536), .clock(clock), .in1(R11535));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11651 (.out1(R11652), .clock(clock), .in1(R11651));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11712 (.out1(R11713), .clock(clock), .in1(R11712));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11768 (.out1(R11769), .clock(clock), .in1(R11768));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11871 (.out1(R11872), .clock(clock), .in1(R11871));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11919 (.out1(R11920), .clock(clock), .in1(R11919));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11962 (.out1(R11963), .clock(clock), .in1(R11962));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12052 (.out1(R12053), .clock(clock), .in1(R12052));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12087 (.out1(R12088), .clock(clock), .in1(R12087));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12117 (.out1(R12118), .clock(clock), .in1(R12117));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12194 (.out1(R12195), .clock(clock), .in1(R12194));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12216 (.out1(R12217), .clock(clock), .in1(R12216));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12233 (.out1(R12234), .clock(clock), .in1(R12233));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12297 (.out1(R12298), .clock(clock), .in1(R12297));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12330 (.out1(R12331), .clock(clock), .in1(_2485));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12331 (.out1(R12332), .clock(clock), .in1(_2390));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12332 (.out1(R12333), .clock(clock), .in1(_2295));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12333 (.out1(R12334), .clock(clock), .in1(_2200));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12334 (.out1(R12335), .clock(clock), .in1(_2105));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12335 (.out1(R12336), .clock(clock), .in1(_2010));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12336 (.out1(R12337), .clock(clock), .in1(_1915));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12337 (.out1(R12338), .clock(clock), .in1(_1820));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12338 (.out1(R12339), .clock(clock), .in1(_1725));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12339 (.out1(R12340), .clock(clock), .in1(_3433));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12340 (.out1(R12341), .clock(clock), .in1(_3338));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12341 (.out1(R12342), .clock(clock), .in1(_1720));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12342 (.out1(R12343), .clock(clock), .in1(_3244));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12343 (.out1(R12344), .clock(clock), .in1(_3149));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12344 (.out1(R12345), .clock(clock), .in1(_3054));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12345 (.out1(R12346), .clock(clock), .in1(_2959));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12346 (.out1(R12347), .clock(clock), .in1(_2864));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12347 (.out1(R12348), .clock(clock), .in1(_2769));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12348 (.out1(R12349), .clock(clock), .in1(_2674));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12349 (.out1(R12350), .clock(clock), .in1(_2579));
  SRAM op3350 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3245),.ADR(R12343));
  SRAM op3252 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3150),.ADR(R12344));
  SRAM op3154 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3055),.ADR(R12345));
  SRAM op3056 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2960),.ADR(R12346));
  SRAM op2958 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2865),.ADR(R12347));
  SRAM op2860 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2770),.ADR(R12348));
  SRAM op2762 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2675),.ADR(R12349));
  SRAM op2664 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2580),.ADR(R12350));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3545 (.out1(_3434), .in1(leafvec16_3539_D), .in2(R12340));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3447 (.out1(_3339), .in1(leafvec22_3548_D), .in2(R12341));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1777 (.out1(_1721), .in1(R12342));
  bit_and #(.BITSIZE_in1(32), .BITSIZE_in2(6), .BITSIZE_out1(32)) op1778 (.out1(off_3683), .in1(_1721), .in2(6 'd 63));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2567 (.out1(_2486), .in1(R12331), .in2(R10494));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2469 (.out1(_2391), .in1(R12332), .in2(R10858));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2371 (.out1(_2296), .in1(R12333), .in2(R11182));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2273 (.out1(_2201), .in1(R12334), .in2(R11467));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2175 (.out1(_2106), .in1(R12335), .in2(R11713));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2077 (.out1(_2011), .in1(R12336), .in2(R11920));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1979 (.out1(_1916), .in1(R12337), .in2(R12088));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1881 (.out1(_1821), .in1(R12338), .in2(R12217));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1783 (.out1(_1726), .in1(R12339), .in2(off_3683));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3928 (.out1(R3929), .clock(clock), .in1(R3928));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4184 (.out1(R4185), .clock(clock), .in1(R4184));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4439 (.out1(R4440), .clock(clock), .in1(R4439));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4684 (.out1(R4685), .clock(clock), .in1(R4684));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4924 (.out1(R4925), .clock(clock), .in1(R4924));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5211 (.out1(R5212), .clock(clock), .in1(R5211));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5443 (.out1(R5444), .clock(clock), .in1(R5443));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5670 (.out1(R5671), .clock(clock), .in1(R5670));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5944 (.out1(R5945), .clock(clock), .in1(R5944));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6162 (.out1(R6163), .clock(clock), .in1(R6162));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6375 (.out1(R6376), .clock(clock), .in1(R6375));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6636 (.out1(R6637), .clock(clock), .in1(R6636));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6841 (.out1(R6842), .clock(clock), .in1(R6841));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7041 (.out1(R7042), .clock(clock), .in1(R7041));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7288 (.out1(R7289), .clock(clock), .in1(R7288));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7480 (.out1(R7481), .clock(clock), .in1(R7480));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7667 (.out1(R7668), .clock(clock), .in1(R7667));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7901 (.out1(R7902), .clock(clock), .in1(R7901));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8080 (.out1(R8081), .clock(clock), .in1(R8080));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8254 (.out1(R8255), .clock(clock), .in1(R8254));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8475 (.out1(R8476), .clock(clock), .in1(R8475));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8641 (.out1(R8642), .clock(clock), .in1(R8641));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8802 (.out1(R8803), .clock(clock), .in1(R8802));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9010 (.out1(R9011), .clock(clock), .in1(R9010));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9163 (.out1(R9164), .clock(clock), .in1(R9163));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9311 (.out1(R9312), .clock(clock), .in1(R9311));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9506 (.out1(R9507), .clock(clock), .in1(R9506));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9646 (.out1(R9647), .clock(clock), .in1(R9646));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9781 (.out1(R9782), .clock(clock), .in1(R9781));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9963 (.out1(R9964), .clock(clock), .in1(R9963));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10090 (.out1(R10091), .clock(clock), .in1(R10090));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10212 (.out1(R10213), .clock(clock), .in1(R10212));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10381 (.out1(R10382), .clock(clock), .in1(R10381));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10494 (.out1(R10495), .clock(clock), .in1(R10494));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10602 (.out1(R10603), .clock(clock), .in1(R10602));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10758 (.out1(R10759), .clock(clock), .in1(R10758));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10858 (.out1(R10859), .clock(clock), .in1(R10858));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10953 (.out1(R10954), .clock(clock), .in1(R10953));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11095 (.out1(R11096), .clock(clock), .in1(R11095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11182 (.out1(R11183), .clock(clock), .in1(R11182));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11264 (.out1(R11265), .clock(clock), .in1(R11264));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11393 (.out1(R11394), .clock(clock), .in1(R11393));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11467 (.out1(R11468), .clock(clock), .in1(R11467));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11536 (.out1(R11537), .clock(clock), .in1(R11536));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11652 (.out1(R11653), .clock(clock), .in1(R11652));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11713 (.out1(R11714), .clock(clock), .in1(R11713));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11769 (.out1(R11770), .clock(clock), .in1(R11769));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11872 (.out1(R11873), .clock(clock), .in1(R11872));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11920 (.out1(R11921), .clock(clock), .in1(R11920));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11963 (.out1(R11964), .clock(clock), .in1(R11963));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12053 (.out1(R12054), .clock(clock), .in1(R12053));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12088 (.out1(R12089), .clock(clock), .in1(R12088));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12118 (.out1(R12119), .clock(clock), .in1(R12118));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12195 (.out1(R12196), .clock(clock), .in1(R12195));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12217 (.out1(R12218), .clock(clock), .in1(R12217));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12234 (.out1(R12235), .clock(clock), .in1(R12234));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12298 (.out1(R12299), .clock(clock), .in1(R12298));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12350 (.out1(R12351), .clock(clock), .in1(_3245));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12351 (.out1(R12352), .clock(clock), .in1(_3150));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12352 (.out1(R12353), .clock(clock), .in1(_3055));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12353 (.out1(R12354), .clock(clock), .in1(_2960));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12354 (.out1(R12355), .clock(clock), .in1(_2865));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12355 (.out1(R12356), .clock(clock), .in1(_2770));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12356 (.out1(R12357), .clock(clock), .in1(_2675));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12357 (.out1(R12358), .clock(clock), .in1(_2580));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12358 (.out1(R12359), .clock(clock), .in1(_3434));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12359 (.out1(R12360), .clock(clock), .in1(_3339));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12360 (.out1(R12361), .clock(clock), .in1(off_3683));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12364 (.out1(R12365), .clock(clock), .in1(_2486));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12365 (.out1(R12366), .clock(clock), .in1(_2391));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12366 (.out1(R12367), .clock(clock), .in1(_2296));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12367 (.out1(R12368), .clock(clock), .in1(_2201));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12368 (.out1(R12369), .clock(clock), .in1(_2106));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12369 (.out1(R12370), .clock(clock), .in1(_2011));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12370 (.out1(R12371), .clock(clock), .in1(_1916));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12371 (.out1(R12372), .clock(clock), .in1(_1821));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12372 (.out1(R12373), .clock(clock), .in1(_1726));
  SRAM op3546 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3435),.ADR(R12359));
  SRAM op3448 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3340),.ADR(R12360));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op2568 (.out1(_2487), .in1(R12365), .in2(1 'd 1));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op2470 (.out1(_2392), .in1(R12366), .in2(1 'd 1));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op2372 (.out1(_2297), .in1(R12367), .in2(1 'd 1));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op2274 (.out1(_2202), .in1(R12368), .in2(1 'd 1));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op2176 (.out1(_2107), .in1(R12369), .in2(1 'd 1));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op2078 (.out1(_2012), .in1(R12370), .in2(1 'd 1));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op1980 (.out1(_1917), .in1(R12371), .in2(1 'd 1));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op1882 (.out1(_1822), .in1(R12372), .in2(1 'd 1));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op1784 (.out1(_1727), .in1(R12373), .in2(1 'd 1));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op2569 (.out1(ifout2569), .in1(_2487), .in2(1 'd 0));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op2471 (.out1(ifout2471), .in1(_2392), .in2(1 'd 0));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op2373 (.out1(ifout2373), .in1(_2297), .in2(1 'd 0));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op2275 (.out1(ifout2275), .in1(_2202), .in2(1 'd 0));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op2177 (.out1(ifout2177), .in1(_2107), .in2(1 'd 0));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op2079 (.out1(ifout2079), .in1(_2012), .in2(1 'd 0));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op1981 (.out1(ifout1981), .in1(_1917), .in2(1 'd 0));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op1883 (.out1(ifout1883), .in1(_1822), .in2(1 'd 0));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op1785 (.out1(ifout1785), .in1(_1727), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2637 (.out1(_2555), .in1(R10382));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2630 (.out1(_2548), .in1(R10382));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2619 (.out1(_2537), .in1(R10382));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2599 (.out1(_2517), .in1(R10382));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2539 (.out1(_2460), .in1(R10759));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2532 (.out1(_2453), .in1(R10759));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2521 (.out1(_2442), .in1(R10759));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2501 (.out1(_2422), .in1(R10759));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2441 (.out1(_2365), .in1(R11096));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2434 (.out1(_2358), .in1(R11096));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2423 (.out1(_2347), .in1(R11096));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2403 (.out1(_2327), .in1(R11096));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2343 (.out1(_2270), .in1(R11394));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2336 (.out1(_2263), .in1(R11394));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2325 (.out1(_2252), .in1(R11394));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2305 (.out1(_2232), .in1(R11394));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2245 (.out1(_2175), .in1(R11653));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2238 (.out1(_2168), .in1(R11653));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2227 (.out1(_2157), .in1(R11653));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2207 (.out1(_2137), .in1(R11653));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2147 (.out1(_2080), .in1(R11873));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2140 (.out1(_2073), .in1(R11873));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2129 (.out1(_2062), .in1(R11873));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2109 (.out1(_2042), .in1(R11873));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2049 (.out1(_1985), .in1(R12054));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2042 (.out1(_1978), .in1(R12054));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2031 (.out1(_1967), .in1(R12054));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2011 (.out1(_1947), .in1(R12054));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1951 (.out1(_1890), .in1(R12196));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1944 (.out1(_1883), .in1(R12196));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1933 (.out1(_1872), .in1(R12196));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1913 (.out1(_1852), .in1(R12196));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1853 (.out1(_1795), .in1(R12299));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1846 (.out1(_1788), .in1(R12299));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1835 (.out1(_1777), .in1(R12299));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1815 (.out1(_1757), .in1(R12299));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2638 (.out1(_2556), .in1(_2555), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2631 (.out1(_2549), .in1(_2548), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2620 (.out1(_2538), .in1(_2537), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2600 (.out1(_2518), .in1(_2517), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2540 (.out1(_2461), .in1(_2460), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2533 (.out1(_2454), .in1(_2453), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2522 (.out1(_2443), .in1(_2442), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2502 (.out1(_2423), .in1(_2422), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2442 (.out1(_2366), .in1(_2365), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2435 (.out1(_2359), .in1(_2358), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2424 (.out1(_2348), .in1(_2347), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2404 (.out1(_2328), .in1(_2327), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2344 (.out1(_2271), .in1(_2270), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2337 (.out1(_2264), .in1(_2263), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2326 (.out1(_2253), .in1(_2252), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2306 (.out1(_2233), .in1(_2232), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2246 (.out1(_2176), .in1(_2175), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2239 (.out1(_2169), .in1(_2168), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2228 (.out1(_2158), .in1(_2157), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2208 (.out1(_2138), .in1(_2137), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2148 (.out1(_2081), .in1(_2080), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2141 (.out1(_2074), .in1(_2073), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2130 (.out1(_2063), .in1(_2062), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2110 (.out1(_2043), .in1(_2042), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2050 (.out1(_1986), .in1(_1985), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2043 (.out1(_1979), .in1(_1978), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2032 (.out1(_1968), .in1(_1967), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2012 (.out1(_1948), .in1(_1947), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1952 (.out1(_1891), .in1(_1890), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1945 (.out1(_1884), .in1(_1883), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1934 (.out1(_1873), .in1(_1872), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1914 (.out1(_1853), .in1(_1852), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1854 (.out1(_1796), .in1(_1795), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1847 (.out1(_1789), .in1(_1788), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1836 (.out1(_1778), .in1(_1777), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1816 (.out1(_1758), .in1(_1757), .in2(2 'd 3));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3351 (.out1(_3246), .in1(R12351), .in2(R6163));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3253 (.out1(_3151), .in1(R12352), .in2(R6842));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3155 (.out1(_3056), .in1(R12353), .in2(R7481));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3057 (.out1(_2961), .in1(R12354), .in2(R8081));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2959 (.out1(_2866), .in1(R12355), .in2(R8642));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2861 (.out1(_2771), .in1(R12356), .in2(R9164));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2763 (.out1(_2676), .in1(R12357), .in2(R9647));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2665 (.out1(_2581), .in1(R12358), .in2(R10091));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3929 (.out1(R3930), .clock(clock), .in1(R3929));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4185 (.out1(R4186), .clock(clock), .in1(R4185));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4440 (.out1(R4441), .clock(clock), .in1(R4440));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4685 (.out1(R4686), .clock(clock), .in1(R4685));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4925 (.out1(R4926), .clock(clock), .in1(R4925));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5212 (.out1(R5213), .clock(clock), .in1(R5212));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5444 (.out1(R5445), .clock(clock), .in1(R5444));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5671 (.out1(R5672), .clock(clock), .in1(R5671));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5945 (.out1(R5946), .clock(clock), .in1(R5945));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6163 (.out1(R6164), .clock(clock), .in1(R6163));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6376 (.out1(R6377), .clock(clock), .in1(R6376));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6637 (.out1(R6638), .clock(clock), .in1(R6637));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6842 (.out1(R6843), .clock(clock), .in1(R6842));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7042 (.out1(R7043), .clock(clock), .in1(R7042));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7289 (.out1(R7290), .clock(clock), .in1(R7289));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7481 (.out1(R7482), .clock(clock), .in1(R7481));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7668 (.out1(R7669), .clock(clock), .in1(R7668));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7902 (.out1(R7903), .clock(clock), .in1(R7902));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8081 (.out1(R8082), .clock(clock), .in1(R8081));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8255 (.out1(R8256), .clock(clock), .in1(R8255));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8476 (.out1(R8477), .clock(clock), .in1(R8476));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8642 (.out1(R8643), .clock(clock), .in1(R8642));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8803 (.out1(R8804), .clock(clock), .in1(R8803));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9011 (.out1(R9012), .clock(clock), .in1(R9011));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9164 (.out1(R9165), .clock(clock), .in1(R9164));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9312 (.out1(R9313), .clock(clock), .in1(R9312));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9507 (.out1(R9508), .clock(clock), .in1(R9507));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9647 (.out1(R9648), .clock(clock), .in1(R9647));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9782 (.out1(R9783), .clock(clock), .in1(R9782));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9964 (.out1(R9965), .clock(clock), .in1(R9964));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10091 (.out1(R10092), .clock(clock), .in1(R10091));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10213 (.out1(R10214), .clock(clock), .in1(R10213));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10382 (.out1(R10383), .clock(clock), .in1(R10382));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10495 (.out1(R10496), .clock(clock), .in1(R10495));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10603 (.out1(R10604), .clock(clock), .in1(R10603));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10759 (.out1(R10760), .clock(clock), .in1(R10759));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10859 (.out1(R10860), .clock(clock), .in1(R10859));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10954 (.out1(R10955), .clock(clock), .in1(R10954));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11096 (.out1(R11097), .clock(clock), .in1(R11096));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11183 (.out1(R11184), .clock(clock), .in1(R11183));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11265 (.out1(R11266), .clock(clock), .in1(R11265));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11394 (.out1(R11395), .clock(clock), .in1(R11394));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11468 (.out1(R11469), .clock(clock), .in1(R11468));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11537 (.out1(R11538), .clock(clock), .in1(R11537));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11653 (.out1(R11654), .clock(clock), .in1(R11653));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11714 (.out1(R11715), .clock(clock), .in1(R11714));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11770 (.out1(R11771), .clock(clock), .in1(R11770));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11873 (.out1(R11874), .clock(clock), .in1(R11873));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11921 (.out1(R11922), .clock(clock), .in1(R11921));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11964 (.out1(R11965), .clock(clock), .in1(R11964));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12054 (.out1(R12055), .clock(clock), .in1(R12054));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12089 (.out1(R12090), .clock(clock), .in1(R12089));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12119 (.out1(R12120), .clock(clock), .in1(R12119));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12196 (.out1(R12197), .clock(clock), .in1(R12196));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12218 (.out1(R12219), .clock(clock), .in1(R12218));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12235 (.out1(R12236), .clock(clock), .in1(R12235));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12299 (.out1(R12300), .clock(clock), .in1(R12299));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12361 (.out1(R12362), .clock(clock), .in1(R12361));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12373 (.out1(R12374), .clock(clock), .in1(_3435));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12374 (.out1(R12375), .clock(clock), .in1(_3340));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12375 (.out1(R12376), .clock(clock), .in1(ifout2569));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12386 (.out1(R12387), .clock(clock), .in1(ifout2471));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12397 (.out1(R12398), .clock(clock), .in1(ifout2373));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12408 (.out1(R12409), .clock(clock), .in1(ifout2275));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12419 (.out1(R12420), .clock(clock), .in1(ifout2177));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12430 (.out1(R12431), .clock(clock), .in1(ifout2079));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12441 (.out1(R12442), .clock(clock), .in1(ifout1981));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12452 (.out1(R12453), .clock(clock), .in1(ifout1883));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12463 (.out1(R12464), .clock(clock), .in1(ifout1785));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12474 (.out1(R12475), .clock(clock), .in1(_2556));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12475 (.out1(R12476), .clock(clock), .in1(_2549));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12476 (.out1(R12477), .clock(clock), .in1(_2538));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12477 (.out1(R12478), .clock(clock), .in1(_2518));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12478 (.out1(R12479), .clock(clock), .in1(_2461));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12479 (.out1(R12480), .clock(clock), .in1(_2454));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12480 (.out1(R12481), .clock(clock), .in1(_2443));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12481 (.out1(R12482), .clock(clock), .in1(_2423));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12482 (.out1(R12483), .clock(clock), .in1(_2366));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12483 (.out1(R12484), .clock(clock), .in1(_2359));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12484 (.out1(R12485), .clock(clock), .in1(_2348));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12485 (.out1(R12486), .clock(clock), .in1(_2328));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12486 (.out1(R12487), .clock(clock), .in1(_2271));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12487 (.out1(R12488), .clock(clock), .in1(_2264));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12488 (.out1(R12489), .clock(clock), .in1(_2253));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12489 (.out1(R12490), .clock(clock), .in1(_2233));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12490 (.out1(R12491), .clock(clock), .in1(_2176));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12491 (.out1(R12492), .clock(clock), .in1(_2169));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12492 (.out1(R12493), .clock(clock), .in1(_2158));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12493 (.out1(R12494), .clock(clock), .in1(_2138));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12494 (.out1(R12495), .clock(clock), .in1(_2081));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12495 (.out1(R12496), .clock(clock), .in1(_2074));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12496 (.out1(R12497), .clock(clock), .in1(_2063));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12497 (.out1(R12498), .clock(clock), .in1(_2043));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12498 (.out1(R12499), .clock(clock), .in1(_1986));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12499 (.out1(R12500), .clock(clock), .in1(_1979));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12500 (.out1(R12501), .clock(clock), .in1(_1968));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12501 (.out1(R12502), .clock(clock), .in1(_1948));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12502 (.out1(R12503), .clock(clock), .in1(_1891));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12503 (.out1(R12504), .clock(clock), .in1(_1884));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12504 (.out1(R12505), .clock(clock), .in1(_1873));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12505 (.out1(R12506), .clock(clock), .in1(_1853));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12506 (.out1(R12507), .clock(clock), .in1(_1796));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12507 (.out1(R12508), .clock(clock), .in1(_1789));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12508 (.out1(R12509), .clock(clock), .in1(_1778));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12509 (.out1(R12510), .clock(clock), .in1(_1758));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12510 (.out1(R12511), .clock(clock), .in1(_3246));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12511 (.out1(R12512), .clock(clock), .in1(_3151));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12512 (.out1(R12513), .clock(clock), .in1(_3056));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12513 (.out1(R12514), .clock(clock), .in1(_2961));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12514 (.out1(R12515), .clock(clock), .in1(_2866));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12515 (.out1(R12516), .clock(clock), .in1(_2771));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12516 (.out1(R12517), .clock(clock), .in1(_2676));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12517 (.out1(R12518), .clock(clock), .in1(_2581));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op3352 (.out1(_3247), .in1(R12511), .in2(1 'd 1));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op3254 (.out1(_3152), .in1(R12512), .in2(1 'd 1));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op3156 (.out1(_3057), .in1(R12513), .in2(1 'd 1));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op3058 (.out1(_2962), .in1(R12514), .in2(1 'd 1));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op2960 (.out1(_2867), .in1(R12515), .in2(1 'd 1));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op2862 (.out1(_2772), .in1(R12516), .in2(1 'd 1));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op2764 (.out1(_2677), .in1(R12517), .in2(1 'd 1));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op2666 (.out1(_2582), .in1(R12518), .in2(1 'd 1));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op3353 (.out1(ifout3353), .in1(_3247), .in2(1 'd 0));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op3255 (.out1(ifout3255), .in1(_3152), .in2(1 'd 0));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op3157 (.out1(ifout3157), .in1(_3057), .in2(1 'd 0));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op3059 (.out1(ifout3059), .in1(_2962), .in2(1 'd 0));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op2961 (.out1(ifout2961), .in1(_2867), .in2(1 'd 0));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op2863 (.out1(ifout2863), .in1(_2772), .in2(1 'd 0));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op2765 (.out1(ifout2765), .in1(_2677), .in2(1 'd 0));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op2667 (.out1(ifout2667), .in1(_2582), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3421 (.out1(_3315), .in1(R5946));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3414 (.out1(_3308), .in1(R5946));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3403 (.out1(_3297), .in1(R5946));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3383 (.out1(_3277), .in1(R5946));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3323 (.out1(_3220), .in1(R6638));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3316 (.out1(_3213), .in1(R6638));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3305 (.out1(_3202), .in1(R6638));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3285 (.out1(_3182), .in1(R6638));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3225 (.out1(_3125), .in1(R7290));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3218 (.out1(_3118), .in1(R7290));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3207 (.out1(_3107), .in1(R7290));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3187 (.out1(_3087), .in1(R7290));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3127 (.out1(_3030), .in1(R7903));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3120 (.out1(_3023), .in1(R7903));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3109 (.out1(_3012), .in1(R7903));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3089 (.out1(_2992), .in1(R7903));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3029 (.out1(_2935), .in1(R8477));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3022 (.out1(_2928), .in1(R8477));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3011 (.out1(_2917), .in1(R8477));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2991 (.out1(_2897), .in1(R8477));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2931 (.out1(_2840), .in1(R9012));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2924 (.out1(_2833), .in1(R9012));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2913 (.out1(_2822), .in1(R9012));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2893 (.out1(_2802), .in1(R9012));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2833 (.out1(_2745), .in1(R9508));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2826 (.out1(_2738), .in1(R9508));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2815 (.out1(_2727), .in1(R9508));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2795 (.out1(_2707), .in1(R9508));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2735 (.out1(_2650), .in1(R9965));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2728 (.out1(_2643), .in1(R9965));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2717 (.out1(_2632), .in1(R9965));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2697 (.out1(_2612), .in1(R9965));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2612 (.out1(_2530), .in1(R10383));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2592 (.out1(_2510), .in1(R10383));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2581 (.out1(_2499), .in1(R10383));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2574 (.out1(_2492), .in1(R10383));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2514 (.out1(_2435), .in1(R10760));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2494 (.out1(_2415), .in1(R10760));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2483 (.out1(_2404), .in1(R10760));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2476 (.out1(_2397), .in1(R10760));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2416 (.out1(_2340), .in1(R11097));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2396 (.out1(_2320), .in1(R11097));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2385 (.out1(_2309), .in1(R11097));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2378 (.out1(_2302), .in1(R11097));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2318 (.out1(_2245), .in1(R11395));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2298 (.out1(_2225), .in1(R11395));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2287 (.out1(_2214), .in1(R11395));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2280 (.out1(_2207), .in1(R11395));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2220 (.out1(_2150), .in1(R11654));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2200 (.out1(_2130), .in1(R11654));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2189 (.out1(_2119), .in1(R11654));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2182 (.out1(_2112), .in1(R11654));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2122 (.out1(_2055), .in1(R11874));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2102 (.out1(_2035), .in1(R11874));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2091 (.out1(_2024), .in1(R11874));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2084 (.out1(_2017), .in1(R11874));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2024 (.out1(_1960), .in1(R12055));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2004 (.out1(_1940), .in1(R12055));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1993 (.out1(_1929), .in1(R12055));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1986 (.out1(_1922), .in1(R12055));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1926 (.out1(_1865), .in1(R12197));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1906 (.out1(_1845), .in1(R12197));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1895 (.out1(_1834), .in1(R12197));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1888 (.out1(_1827), .in1(R12197));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1828 (.out1(_1770), .in1(R12300));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1808 (.out1(_1750), .in1(R12300));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1797 (.out1(_1739), .in1(R12300));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1790 (.out1(_1732), .in1(R12300));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3422 (.out1(_3316), .in1(_3315), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3415 (.out1(_3309), .in1(_3308), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3404 (.out1(_3298), .in1(_3297), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3384 (.out1(_3278), .in1(_3277), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3324 (.out1(_3221), .in1(_3220), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3317 (.out1(_3214), .in1(_3213), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3306 (.out1(_3203), .in1(_3202), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3286 (.out1(_3183), .in1(_3182), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3226 (.out1(_3126), .in1(_3125), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3219 (.out1(_3119), .in1(_3118), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3208 (.out1(_3108), .in1(_3107), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3188 (.out1(_3088), .in1(_3087), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3128 (.out1(_3031), .in1(_3030), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3121 (.out1(_3024), .in1(_3023), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3110 (.out1(_3013), .in1(_3012), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3090 (.out1(_2993), .in1(_2992), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3030 (.out1(_2936), .in1(_2935), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3023 (.out1(_2929), .in1(_2928), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3012 (.out1(_2918), .in1(_2917), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2992 (.out1(_2898), .in1(_2897), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2932 (.out1(_2841), .in1(_2840), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2925 (.out1(_2834), .in1(_2833), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2914 (.out1(_2823), .in1(_2822), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2894 (.out1(_2803), .in1(_2802), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2834 (.out1(_2746), .in1(_2745), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2827 (.out1(_2739), .in1(_2738), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2816 (.out1(_2728), .in1(_2727), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2796 (.out1(_2708), .in1(_2707), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2736 (.out1(_2651), .in1(_2650), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2729 (.out1(_2644), .in1(_2643), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2718 (.out1(_2633), .in1(_2632), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2698 (.out1(_2613), .in1(_2612), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2641 (.out1(_2559), .in1(2 'd 2), .in2(R10496));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2613 (.out1(_2531), .in1(_2530), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2593 (.out1(_2511), .in1(_2510), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2582 (.out1(_2500), .in1(_2499), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2575 (.out1(_2493), .in1(_2492), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2543 (.out1(_2464), .in1(2 'd 2), .in2(R10860));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2515 (.out1(_2436), .in1(_2435), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2495 (.out1(_2416), .in1(_2415), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2484 (.out1(_2405), .in1(_2404), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2477 (.out1(_2398), .in1(_2397), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2445 (.out1(_2369), .in1(2 'd 2), .in2(R11184));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2417 (.out1(_2341), .in1(_2340), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2397 (.out1(_2321), .in1(_2320), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2386 (.out1(_2310), .in1(_2309), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2379 (.out1(_2303), .in1(_2302), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2347 (.out1(_2274), .in1(2 'd 2), .in2(R11469));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2319 (.out1(_2246), .in1(_2245), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2299 (.out1(_2226), .in1(_2225), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2288 (.out1(_2215), .in1(_2214), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2281 (.out1(_2208), .in1(_2207), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2249 (.out1(_2179), .in1(2 'd 2), .in2(R11715));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2221 (.out1(_2151), .in1(_2150), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2201 (.out1(_2131), .in1(_2130), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2190 (.out1(_2120), .in1(_2119), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2183 (.out1(_2113), .in1(_2112), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2151 (.out1(_2084), .in1(2 'd 2), .in2(R11922));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2123 (.out1(_2056), .in1(_2055), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2103 (.out1(_2036), .in1(_2035), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2092 (.out1(_2025), .in1(_2024), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2085 (.out1(_2018), .in1(_2017), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2053 (.out1(_1989), .in1(2 'd 2), .in2(R12090));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2025 (.out1(_1961), .in1(_1960), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2005 (.out1(_1941), .in1(_1940), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1994 (.out1(_1930), .in1(_1929), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1987 (.out1(_1923), .in1(_1922), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1955 (.out1(_1894), .in1(2 'd 2), .in2(R12219));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1927 (.out1(_1866), .in1(_1865), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1907 (.out1(_1846), .in1(_1845), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1896 (.out1(_1835), .in1(_1834), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1889 (.out1(_1828), .in1(_1827), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1857 (.out1(_1799), .in1(2 'd 2), .in2(R12362));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1829 (.out1(_1771), .in1(_1770), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1809 (.out1(_1751), .in1(_1750), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1798 (.out1(_1740), .in1(_1739), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1791 (.out1(_1733), .in1(_1732), .in2(2 'd 3));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2639 (.out1(_2557), .in1(leafvec76_3621_D), .in2(R12475));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2632 (.out1(_2550), .in1(leafvec76_3621_D), .in2(R12476));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2621 (.out1(_2539), .in1(leafvec76_3621_D), .in2(R12477));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2601 (.out1(_2519), .in1(leafvec76_3621_D), .in2(R12478));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2541 (.out1(_2462), .in1(leafvec82_3629_D), .in2(R12479));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2534 (.out1(_2455), .in1(leafvec82_3629_D), .in2(R12480));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2523 (.out1(_2444), .in1(leafvec82_3629_D), .in2(R12481));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2503 (.out1(_2424), .in1(leafvec82_3629_D), .in2(R12482));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2443 (.out1(_2367), .in1(leafvec88_3637_D), .in2(R12483));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2436 (.out1(_2360), .in1(leafvec88_3637_D), .in2(R12484));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2425 (.out1(_2349), .in1(leafvec88_3637_D), .in2(R12485));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2405 (.out1(_2329), .in1(leafvec88_3637_D), .in2(R12486));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2345 (.out1(_2272), .in1(leafvec94_3645_D), .in2(R12487));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2338 (.out1(_2265), .in1(leafvec94_3645_D), .in2(R12488));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2327 (.out1(_2254), .in1(leafvec94_3645_D), .in2(R12489));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2307 (.out1(_2234), .in1(leafvec94_3645_D), .in2(R12490));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2247 (.out1(_2177), .in1(leafvec100_3653_D), .in2(R12491));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2240 (.out1(_2170), .in1(leafvec100_3653_D), .in2(R12492));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2229 (.out1(_2159), .in1(leafvec100_3653_D), .in2(R12493));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2209 (.out1(_2139), .in1(leafvec100_3653_D), .in2(R12494));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2149 (.out1(_2082), .in1(leafvec106_3661_D), .in2(R12495));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2142 (.out1(_2075), .in1(leafvec106_3661_D), .in2(R12496));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2131 (.out1(_2064), .in1(leafvec106_3661_D), .in2(R12497));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2111 (.out1(_2044), .in1(leafvec106_3661_D), .in2(R12498));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2051 (.out1(_1987), .in1(leafvec112_3669_D), .in2(R12499));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2044 (.out1(_1980), .in1(leafvec112_3669_D), .in2(R12500));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2033 (.out1(_1969), .in1(leafvec112_3669_D), .in2(R12501));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2013 (.out1(_1949), .in1(leafvec112_3669_D), .in2(R12502));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1953 (.out1(_1892), .in1(leafvec118_3677_D), .in2(R12503));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1946 (.out1(_1885), .in1(leafvec118_3677_D), .in2(R12504));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1935 (.out1(_1874), .in1(leafvec118_3677_D), .in2(R12505));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1915 (.out1(_1854), .in1(leafvec118_3677_D), .in2(R12506));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1855 (.out1(_1797), .in1(leafvec124_3684_D), .in2(R12507));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1848 (.out1(_1790), .in1(leafvec124_3684_D), .in2(R12508));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1837 (.out1(_1779), .in1(leafvec124_3684_D), .in2(R12509));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1817 (.out1(_1759), .in1(leafvec124_3684_D), .in2(R12510));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3547 (.out1(_3436), .in1(R12374), .in2(R4686));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3449 (.out1(_3341), .in1(R12375), .in2(R5445));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3930 (.out1(R3931), .clock(clock), .in1(R3930));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4186 (.out1(R4187), .clock(clock), .in1(R4186));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4441 (.out1(R4442), .clock(clock), .in1(R4441));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4686 (.out1(R4687), .clock(clock), .in1(R4686));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4926 (.out1(R4927), .clock(clock), .in1(R4926));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5213 (.out1(R5214), .clock(clock), .in1(R5213));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5445 (.out1(R5446), .clock(clock), .in1(R5445));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5672 (.out1(R5673), .clock(clock), .in1(R5672));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5946 (.out1(R5947), .clock(clock), .in1(R5946));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6164 (.out1(R6165), .clock(clock), .in1(R6164));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6377 (.out1(R6378), .clock(clock), .in1(R6377));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6638 (.out1(R6639), .clock(clock), .in1(R6638));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6843 (.out1(R6844), .clock(clock), .in1(R6843));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7043 (.out1(R7044), .clock(clock), .in1(R7043));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7290 (.out1(R7291), .clock(clock), .in1(R7290));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7482 (.out1(R7483), .clock(clock), .in1(R7482));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7669 (.out1(R7670), .clock(clock), .in1(R7669));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7903 (.out1(R7904), .clock(clock), .in1(R7903));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8082 (.out1(R8083), .clock(clock), .in1(R8082));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8256 (.out1(R8257), .clock(clock), .in1(R8256));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8477 (.out1(R8478), .clock(clock), .in1(R8477));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8643 (.out1(R8644), .clock(clock), .in1(R8643));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8804 (.out1(R8805), .clock(clock), .in1(R8804));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9012 (.out1(R9013), .clock(clock), .in1(R9012));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9165 (.out1(R9166), .clock(clock), .in1(R9165));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9313 (.out1(R9314), .clock(clock), .in1(R9313));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9508 (.out1(R9509), .clock(clock), .in1(R9508));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9648 (.out1(R9649), .clock(clock), .in1(R9648));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9783 (.out1(R9784), .clock(clock), .in1(R9783));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9965 (.out1(R9966), .clock(clock), .in1(R9965));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10092 (.out1(R10093), .clock(clock), .in1(R10092));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10214 (.out1(R10215), .clock(clock), .in1(R10214));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10383 (.out1(R10384), .clock(clock), .in1(R10383));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10496 (.out1(R10497), .clock(clock), .in1(R10496));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10604 (.out1(R10605), .clock(clock), .in1(R10604));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10760 (.out1(R10761), .clock(clock), .in1(R10760));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10860 (.out1(R10861), .clock(clock), .in1(R10860));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10955 (.out1(R10956), .clock(clock), .in1(R10955));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11097 (.out1(R11098), .clock(clock), .in1(R11097));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11184 (.out1(R11185), .clock(clock), .in1(R11184));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11266 (.out1(R11267), .clock(clock), .in1(R11266));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11395 (.out1(R11396), .clock(clock), .in1(R11395));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11469 (.out1(R11470), .clock(clock), .in1(R11469));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11538 (.out1(R11539), .clock(clock), .in1(R11538));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11654 (.out1(R11655), .clock(clock), .in1(R11654));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11715 (.out1(R11716), .clock(clock), .in1(R11715));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11771 (.out1(R11772), .clock(clock), .in1(R11771));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11874 (.out1(R11875), .clock(clock), .in1(R11874));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11922 (.out1(R11923), .clock(clock), .in1(R11922));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11965 (.out1(R11966), .clock(clock), .in1(R11965));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12055 (.out1(R12056), .clock(clock), .in1(R12055));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12090 (.out1(R12091), .clock(clock), .in1(R12090));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12120 (.out1(R12121), .clock(clock), .in1(R12120));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12197 (.out1(R12198), .clock(clock), .in1(R12197));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12219 (.out1(R12220), .clock(clock), .in1(R12219));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12236 (.out1(R12237), .clock(clock), .in1(R12236));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12300 (.out1(R12301), .clock(clock), .in1(R12300));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12362 (.out1(R12363), .clock(clock), .in1(R12362));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12376 (.out1(R12377), .clock(clock), .in1(R12376));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12387 (.out1(R12388), .clock(clock), .in1(R12387));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12398 (.out1(R12399), .clock(clock), .in1(R12398));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12409 (.out1(R12410), .clock(clock), .in1(R12409));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12420 (.out1(R12421), .clock(clock), .in1(R12420));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12431 (.out1(R12432), .clock(clock), .in1(R12431));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12442 (.out1(R12443), .clock(clock), .in1(R12442));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12453 (.out1(R12454), .clock(clock), .in1(R12453));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12464 (.out1(R12465), .clock(clock), .in1(R12464));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12518 (.out1(R12519), .clock(clock), .in1(ifout3353));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12529 (.out1(R12530), .clock(clock), .in1(ifout3255));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12540 (.out1(R12541), .clock(clock), .in1(ifout3157));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12551 (.out1(R12552), .clock(clock), .in1(ifout3059));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12562 (.out1(R12563), .clock(clock), .in1(ifout2961));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12573 (.out1(R12574), .clock(clock), .in1(ifout2863));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12584 (.out1(R12585), .clock(clock), .in1(ifout2765));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12595 (.out1(R12596), .clock(clock), .in1(ifout2667));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12606 (.out1(R12607), .clock(clock), .in1(_3316));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12607 (.out1(R12608), .clock(clock), .in1(_3309));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12608 (.out1(R12609), .clock(clock), .in1(_3298));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12609 (.out1(R12610), .clock(clock), .in1(_3278));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12610 (.out1(R12611), .clock(clock), .in1(_3221));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12611 (.out1(R12612), .clock(clock), .in1(_3214));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12612 (.out1(R12613), .clock(clock), .in1(_3203));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12613 (.out1(R12614), .clock(clock), .in1(_3183));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12614 (.out1(R12615), .clock(clock), .in1(_3126));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12615 (.out1(R12616), .clock(clock), .in1(_3119));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12616 (.out1(R12617), .clock(clock), .in1(_3108));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12617 (.out1(R12618), .clock(clock), .in1(_3088));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12618 (.out1(R12619), .clock(clock), .in1(_3031));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12619 (.out1(R12620), .clock(clock), .in1(_3024));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12620 (.out1(R12621), .clock(clock), .in1(_3013));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12621 (.out1(R12622), .clock(clock), .in1(_2993));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12622 (.out1(R12623), .clock(clock), .in1(_2936));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12623 (.out1(R12624), .clock(clock), .in1(_2929));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12624 (.out1(R12625), .clock(clock), .in1(_2918));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12625 (.out1(R12626), .clock(clock), .in1(_2898));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12626 (.out1(R12627), .clock(clock), .in1(_2841));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12627 (.out1(R12628), .clock(clock), .in1(_2834));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12628 (.out1(R12629), .clock(clock), .in1(_2823));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12629 (.out1(R12630), .clock(clock), .in1(_2803));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12630 (.out1(R12631), .clock(clock), .in1(_2746));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12631 (.out1(R12632), .clock(clock), .in1(_2739));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12632 (.out1(R12633), .clock(clock), .in1(_2728));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12633 (.out1(R12634), .clock(clock), .in1(_2708));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12634 (.out1(R12635), .clock(clock), .in1(_2651));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12635 (.out1(R12636), .clock(clock), .in1(_2644));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12636 (.out1(R12637), .clock(clock), .in1(_2633));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12637 (.out1(R12638), .clock(clock), .in1(_2613));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12638 (.out1(R12639), .clock(clock), .in1(_2559));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12639 (.out1(R12640), .clock(clock), .in1(_2531));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12640 (.out1(R12641), .clock(clock), .in1(_2511));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12641 (.out1(R12642), .clock(clock), .in1(_2500));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12642 (.out1(R12643), .clock(clock), .in1(_2493));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12643 (.out1(R12644), .clock(clock), .in1(_2464));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12644 (.out1(R12645), .clock(clock), .in1(_2436));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12645 (.out1(R12646), .clock(clock), .in1(_2416));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12646 (.out1(R12647), .clock(clock), .in1(_2405));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12647 (.out1(R12648), .clock(clock), .in1(_2398));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12648 (.out1(R12649), .clock(clock), .in1(_2369));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12649 (.out1(R12650), .clock(clock), .in1(_2341));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12650 (.out1(R12651), .clock(clock), .in1(_2321));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12651 (.out1(R12652), .clock(clock), .in1(_2310));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12652 (.out1(R12653), .clock(clock), .in1(_2303));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12653 (.out1(R12654), .clock(clock), .in1(_2274));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12654 (.out1(R12655), .clock(clock), .in1(_2246));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12655 (.out1(R12656), .clock(clock), .in1(_2226));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12656 (.out1(R12657), .clock(clock), .in1(_2215));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12657 (.out1(R12658), .clock(clock), .in1(_2208));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12658 (.out1(R12659), .clock(clock), .in1(_2179));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12659 (.out1(R12660), .clock(clock), .in1(_2151));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12660 (.out1(R12661), .clock(clock), .in1(_2131));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12661 (.out1(R12662), .clock(clock), .in1(_2120));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12662 (.out1(R12663), .clock(clock), .in1(_2113));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12663 (.out1(R12664), .clock(clock), .in1(_2084));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12664 (.out1(R12665), .clock(clock), .in1(_2056));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12665 (.out1(R12666), .clock(clock), .in1(_2036));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12666 (.out1(R12667), .clock(clock), .in1(_2025));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12667 (.out1(R12668), .clock(clock), .in1(_2018));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12668 (.out1(R12669), .clock(clock), .in1(_1989));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12669 (.out1(R12670), .clock(clock), .in1(_1961));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12670 (.out1(R12671), .clock(clock), .in1(_1941));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12671 (.out1(R12672), .clock(clock), .in1(_1930));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12672 (.out1(R12673), .clock(clock), .in1(_1923));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12673 (.out1(R12674), .clock(clock), .in1(_1894));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12674 (.out1(R12675), .clock(clock), .in1(_1866));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12675 (.out1(R12676), .clock(clock), .in1(_1846));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12676 (.out1(R12677), .clock(clock), .in1(_1835));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12677 (.out1(R12678), .clock(clock), .in1(_1828));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12678 (.out1(R12679), .clock(clock), .in1(_1799));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12679 (.out1(R12680), .clock(clock), .in1(_1771));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12680 (.out1(R12681), .clock(clock), .in1(_1751));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12681 (.out1(R12682), .clock(clock), .in1(_1740));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12682 (.out1(R12683), .clock(clock), .in1(_1733));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12683 (.out1(R12684), .clock(clock), .in1(_2557));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12684 (.out1(R12685), .clock(clock), .in1(_2550));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12685 (.out1(R12686), .clock(clock), .in1(_2539));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12686 (.out1(R12687), .clock(clock), .in1(_2519));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12687 (.out1(R12688), .clock(clock), .in1(_2462));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12688 (.out1(R12689), .clock(clock), .in1(_2455));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12689 (.out1(R12690), .clock(clock), .in1(_2444));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12690 (.out1(R12691), .clock(clock), .in1(_2424));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12691 (.out1(R12692), .clock(clock), .in1(_2367));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12692 (.out1(R12693), .clock(clock), .in1(_2360));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12693 (.out1(R12694), .clock(clock), .in1(_2349));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12694 (.out1(R12695), .clock(clock), .in1(_2329));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12695 (.out1(R12696), .clock(clock), .in1(_2272));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12696 (.out1(R12697), .clock(clock), .in1(_2265));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12697 (.out1(R12698), .clock(clock), .in1(_2254));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12698 (.out1(R12699), .clock(clock), .in1(_2234));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12699 (.out1(R12700), .clock(clock), .in1(_2177));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12700 (.out1(R12701), .clock(clock), .in1(_2170));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12701 (.out1(R12702), .clock(clock), .in1(_2159));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12702 (.out1(R12703), .clock(clock), .in1(_2139));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12703 (.out1(R12704), .clock(clock), .in1(_2082));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12704 (.out1(R12705), .clock(clock), .in1(_2075));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12705 (.out1(R12706), .clock(clock), .in1(_2064));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12706 (.out1(R12707), .clock(clock), .in1(_2044));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12707 (.out1(R12708), .clock(clock), .in1(_1987));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12708 (.out1(R12709), .clock(clock), .in1(_1980));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12709 (.out1(R12710), .clock(clock), .in1(_1969));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12710 (.out1(R12711), .clock(clock), .in1(_1949));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12711 (.out1(R12712), .clock(clock), .in1(_1892));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12712 (.out1(R12713), .clock(clock), .in1(_1885));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12713 (.out1(R12714), .clock(clock), .in1(_1874));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12714 (.out1(R12715), .clock(clock), .in1(_1854));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12715 (.out1(R12716), .clock(clock), .in1(_1797));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12716 (.out1(R12717), .clock(clock), .in1(_1790));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12717 (.out1(R12718), .clock(clock), .in1(_1779));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12718 (.out1(R12719), .clock(clock), .in1(_1759));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12719 (.out1(R12720), .clock(clock), .in1(_3436));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12720 (.out1(R12721), .clock(clock), .in1(_3341));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op3548 (.out1(_3437), .in1(R12720), .in2(1 'd 1));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64)) op3450 (.out1(_3342), .in1(R12721), .in2(1 'd 1));
  SRAM op2640 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2558),.ADR(R12684));
  SRAM op2633 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2551),.ADR(R12685));
  SRAM op2622 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2540),.ADR(R12686));
  SRAM op2602 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2520),.ADR(R12687));
  SRAM op2542 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2463),.ADR(R12688));
  SRAM op2535 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2456),.ADR(R12689));
  SRAM op2524 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2445),.ADR(R12690));
  SRAM op2504 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2425),.ADR(R12691));
  SRAM op2444 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2368),.ADR(R12692));
  SRAM op2437 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2361),.ADR(R12693));
  SRAM op2426 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2350),.ADR(R12694));
  SRAM op2406 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2330),.ADR(R12695));
  SRAM op2346 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2273),.ADR(R12696));
  SRAM op2339 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2266),.ADR(R12697));
  SRAM op2328 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2255),.ADR(R12698));
  SRAM op2308 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2235),.ADR(R12699));
  SRAM op2248 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2178),.ADR(R12700));
  SRAM op2241 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2171),.ADR(R12701));
  SRAM op2230 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2160),.ADR(R12702));
  SRAM op2210 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2140),.ADR(R12703));
  SRAM op2150 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2083),.ADR(R12704));
  SRAM op2143 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2076),.ADR(R12705));
  SRAM op2132 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2065),.ADR(R12706));
  SRAM op2112 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2045),.ADR(R12707));
  SRAM op2052 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1988),.ADR(R12708));
  SRAM op2045 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1981),.ADR(R12709));
  SRAM op2034 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1970),.ADR(R12710));
  SRAM op2014 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1950),.ADR(R12711));
  SRAM op1954 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1893),.ADR(R12712));
  SRAM op1947 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1886),.ADR(R12713));
  SRAM op1936 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1875),.ADR(R12714));
  SRAM op1916 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1855),.ADR(R12715));
  SRAM op1856 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1798),.ADR(R12716));
  SRAM op1849 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1791),.ADR(R12717));
  SRAM op1838 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1780),.ADR(R12718));
  SRAM op1818 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1760),.ADR(R12719));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op3549 (.out1(ifout3549), .in1(_3437), .in2(1 'd 0));
  NE_EXPR #(.BITSIZE_in1(64), .BITSIZE_in2(1),.BITSIZE_out1(1)) op3451 (.out1(ifout3451), .in1(_3342), .in2(1 'd 0));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3617 (.out1(_3505), .in1(R4442));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3610 (.out1(_3498), .in1(R4442));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3599 (.out1(_3487), .in1(R4442));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3579 (.out1(_3467), .in1(R4442));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3519 (.out1(_3410), .in1(R5214));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3512 (.out1(_3403), .in1(R5214));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3501 (.out1(_3392), .in1(R5214));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3481 (.out1(_3372), .in1(R5214));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3396 (.out1(_3290), .in1(R5947));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3376 (.out1(_3270), .in1(R5947));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3365 (.out1(_3259), .in1(R5947));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3358 (.out1(_3252), .in1(R5947));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3298 (.out1(_3195), .in1(R6639));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3278 (.out1(_3175), .in1(R6639));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3267 (.out1(_3164), .in1(R6639));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3260 (.out1(_3157), .in1(R6639));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3200 (.out1(_3100), .in1(R7291));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3180 (.out1(_3080), .in1(R7291));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3169 (.out1(_3069), .in1(R7291));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3162 (.out1(_3062), .in1(R7291));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3102 (.out1(_3005), .in1(R7904));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3082 (.out1(_2985), .in1(R7904));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3071 (.out1(_2974), .in1(R7904));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3064 (.out1(_2967), .in1(R7904));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3004 (.out1(_2910), .in1(R8478));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2984 (.out1(_2890), .in1(R8478));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2973 (.out1(_2879), .in1(R8478));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2966 (.out1(_2872), .in1(R8478));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2906 (.out1(_2815), .in1(R9013));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2886 (.out1(_2795), .in1(R9013));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2875 (.out1(_2784), .in1(R9013));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2868 (.out1(_2777), .in1(R9013));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2808 (.out1(_2720), .in1(R9509));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2788 (.out1(_2700), .in1(R9509));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2777 (.out1(_2689), .in1(R9509));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2770 (.out1(_2682), .in1(R9509));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2710 (.out1(_2625), .in1(R9966));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2690 (.out1(_2605), .in1(R9966));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2679 (.out1(_2594), .in1(R9966));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2672 (.out1(_2587), .in1(R9966));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3618 (.out1(_3506), .in1(_3505), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3611 (.out1(_3499), .in1(_3498), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3600 (.out1(_3488), .in1(_3487), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3580 (.out1(_3468), .in1(_3467), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3520 (.out1(_3411), .in1(_3410), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3513 (.out1(_3404), .in1(_3403), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3502 (.out1(_3393), .in1(_3392), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3482 (.out1(_3373), .in1(_3372), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3425 (.out1(_3319), .in1(2 'd 2), .in2(R6165));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3397 (.out1(_3291), .in1(_3290), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3377 (.out1(_3271), .in1(_3270), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3366 (.out1(_3260), .in1(_3259), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3359 (.out1(_3253), .in1(_3252), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3327 (.out1(_3224), .in1(2 'd 2), .in2(R6844));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3299 (.out1(_3196), .in1(_3195), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3279 (.out1(_3176), .in1(_3175), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3268 (.out1(_3165), .in1(_3164), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3261 (.out1(_3158), .in1(_3157), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3229 (.out1(_3129), .in1(2 'd 2), .in2(R7483));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3201 (.out1(_3101), .in1(_3100), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3181 (.out1(_3081), .in1(_3080), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3170 (.out1(_3070), .in1(_3069), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3163 (.out1(_3063), .in1(_3062), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3131 (.out1(_3034), .in1(2 'd 2), .in2(R8083));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3103 (.out1(_3006), .in1(_3005), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3083 (.out1(_2986), .in1(_2985), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3072 (.out1(_2975), .in1(_2974), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3065 (.out1(_2968), .in1(_2967), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3033 (.out1(_2939), .in1(2 'd 2), .in2(R8644));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3005 (.out1(_2911), .in1(_2910), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2985 (.out1(_2891), .in1(_2890), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2974 (.out1(_2880), .in1(_2879), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2967 (.out1(_2873), .in1(_2872), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2935 (.out1(_2844), .in1(2 'd 2), .in2(R9166));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2907 (.out1(_2816), .in1(_2815), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2887 (.out1(_2796), .in1(_2795), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2876 (.out1(_2785), .in1(_2784), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2869 (.out1(_2778), .in1(_2777), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2837 (.out1(_2749), .in1(2 'd 2), .in2(R9649));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2809 (.out1(_2721), .in1(_2720), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2789 (.out1(_2701), .in1(_2700), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2778 (.out1(_2690), .in1(_2689), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2771 (.out1(_2683), .in1(_2682), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2739 (.out1(_2654), .in1(2 'd 2), .in2(R10093));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2711 (.out1(_2626), .in1(_2625), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2691 (.out1(_2606), .in1(_2605), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2680 (.out1(_2595), .in1(_2594), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2673 (.out1(_2588), .in1(_2587), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2634 (.out1(_2552), .in1(2 'd 2), .in2(R10497));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2623 (.out1(_2541), .in1(2 'd 2), .in2(R10497));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2616 (.out1(_2534), .in1(2 'd 2), .in2(R10497));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2603 (.out1(_2521), .in1(2 'd 2), .in2(R10497));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2596 (.out1(_2514), .in1(2 'd 2), .in2(R10497));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2585 (.out1(_2503), .in1(2 'd 2), .in2(R10497));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2536 (.out1(_2457), .in1(2 'd 2), .in2(R10861));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2525 (.out1(_2446), .in1(2 'd 2), .in2(R10861));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2518 (.out1(_2439), .in1(2 'd 2), .in2(R10861));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2505 (.out1(_2426), .in1(2 'd 2), .in2(R10861));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2498 (.out1(_2419), .in1(2 'd 2), .in2(R10861));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2487 (.out1(_2408), .in1(2 'd 2), .in2(R10861));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2438 (.out1(_2362), .in1(2 'd 2), .in2(R11185));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2427 (.out1(_2351), .in1(2 'd 2), .in2(R11185));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2420 (.out1(_2344), .in1(2 'd 2), .in2(R11185));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2407 (.out1(_2331), .in1(2 'd 2), .in2(R11185));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2400 (.out1(_2324), .in1(2 'd 2), .in2(R11185));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2389 (.out1(_2313), .in1(2 'd 2), .in2(R11185));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2340 (.out1(_2267), .in1(2 'd 2), .in2(R11470));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2329 (.out1(_2256), .in1(2 'd 2), .in2(R11470));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2322 (.out1(_2249), .in1(2 'd 2), .in2(R11470));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2309 (.out1(_2236), .in1(2 'd 2), .in2(R11470));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2302 (.out1(_2229), .in1(2 'd 2), .in2(R11470));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2291 (.out1(_2218), .in1(2 'd 2), .in2(R11470));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2242 (.out1(_2172), .in1(2 'd 2), .in2(R11716));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2231 (.out1(_2161), .in1(2 'd 2), .in2(R11716));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2224 (.out1(_2154), .in1(2 'd 2), .in2(R11716));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2211 (.out1(_2141), .in1(2 'd 2), .in2(R11716));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2204 (.out1(_2134), .in1(2 'd 2), .in2(R11716));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2193 (.out1(_2123), .in1(2 'd 2), .in2(R11716));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2144 (.out1(_2077), .in1(2 'd 2), .in2(R11923));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2133 (.out1(_2066), .in1(2 'd 2), .in2(R11923));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2126 (.out1(_2059), .in1(2 'd 2), .in2(R11923));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2113 (.out1(_2046), .in1(2 'd 2), .in2(R11923));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2106 (.out1(_2039), .in1(2 'd 2), .in2(R11923));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2095 (.out1(_2028), .in1(2 'd 2), .in2(R11923));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2046 (.out1(_1982), .in1(2 'd 2), .in2(R12091));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2035 (.out1(_1971), .in1(2 'd 2), .in2(R12091));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2028 (.out1(_1964), .in1(2 'd 2), .in2(R12091));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2015 (.out1(_1951), .in1(2 'd 2), .in2(R12091));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2008 (.out1(_1944), .in1(2 'd 2), .in2(R12091));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1997 (.out1(_1933), .in1(2 'd 2), .in2(R12091));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1948 (.out1(_1887), .in1(2 'd 2), .in2(R12220));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1937 (.out1(_1876), .in1(2 'd 2), .in2(R12220));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1930 (.out1(_1869), .in1(2 'd 2), .in2(R12220));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1917 (.out1(_1856), .in1(2 'd 2), .in2(R12220));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1910 (.out1(_1849), .in1(2 'd 2), .in2(R12220));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1899 (.out1(_1838), .in1(2 'd 2), .in2(R12220));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1850 (.out1(_1792), .in1(2 'd 2), .in2(R12363));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1839 (.out1(_1781), .in1(2 'd 2), .in2(R12363));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1832 (.out1(_1774), .in1(2 'd 2), .in2(R12363));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1819 (.out1(_1761), .in1(2 'd 2), .in2(R12363));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1812 (.out1(_1754), .in1(2 'd 2), .in2(R12363));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1801 (.out1(_1743), .in1(2 'd 2), .in2(R12363));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3423 (.out1(_3317), .in1(leafvec28_3556_D), .in2(R12607));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3416 (.out1(_3310), .in1(leafvec28_3556_D), .in2(R12608));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3405 (.out1(_3299), .in1(leafvec28_3556_D), .in2(R12609));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3385 (.out1(_3279), .in1(leafvec28_3556_D), .in2(R12610));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3325 (.out1(_3222), .in1(leafvec34_3564_D), .in2(R12611));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3318 (.out1(_3215), .in1(leafvec34_3564_D), .in2(R12612));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3307 (.out1(_3204), .in1(leafvec34_3564_D), .in2(R12613));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3287 (.out1(_3184), .in1(leafvec34_3564_D), .in2(R12614));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3227 (.out1(_3127), .in1(leafvec40_3572_D), .in2(R12615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3220 (.out1(_3120), .in1(leafvec40_3572_D), .in2(R12616));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3209 (.out1(_3109), .in1(leafvec40_3572_D), .in2(R12617));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3189 (.out1(_3089), .in1(leafvec40_3572_D), .in2(R12618));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3129 (.out1(_3032), .in1(leafvec46_3580_D), .in2(R12619));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3122 (.out1(_3025), .in1(leafvec46_3580_D), .in2(R12620));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3111 (.out1(_3014), .in1(leafvec46_3580_D), .in2(R12621));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3091 (.out1(_2994), .in1(leafvec46_3580_D), .in2(R12622));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3031 (.out1(_2937), .in1(leafvec52_3588_D), .in2(R12623));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3024 (.out1(_2930), .in1(leafvec52_3588_D), .in2(R12624));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3013 (.out1(_2919), .in1(leafvec52_3588_D), .in2(R12625));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2993 (.out1(_2899), .in1(leafvec52_3588_D), .in2(R12626));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2933 (.out1(_2842), .in1(leafvec58_3596_D), .in2(R12627));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2926 (.out1(_2835), .in1(leafvec58_3596_D), .in2(R12628));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2915 (.out1(_2824), .in1(leafvec58_3596_D), .in2(R12629));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2895 (.out1(_2804), .in1(leafvec58_3596_D), .in2(R12630));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2835 (.out1(_2747), .in1(leafvec64_3605_D), .in2(R12631));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2828 (.out1(_2740), .in1(leafvec64_3605_D), .in2(R12632));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2817 (.out1(_2729), .in1(leafvec64_3605_D), .in2(R12633));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2797 (.out1(_2709), .in1(leafvec64_3605_D), .in2(R12634));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2737 (.out1(_2652), .in1(leafvec70_3613_D), .in2(R12635));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2730 (.out1(_2645), .in1(leafvec70_3613_D), .in2(R12636));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2719 (.out1(_2634), .in1(leafvec70_3613_D), .in2(R12637));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2699 (.out1(_2614), .in1(leafvec70_3613_D), .in2(R12638));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2614 (.out1(_2532), .in1(leafvec76_3621_D), .in2(R12640));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2594 (.out1(_2512), .in1(leafvec76_3621_D), .in2(R12641));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2583 (.out1(_2501), .in1(leafvec76_3621_D), .in2(R12642));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2576 (.out1(_2494), .in1(leafvec76_3621_D), .in2(R12643));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2516 (.out1(_2437), .in1(leafvec82_3629_D), .in2(R12645));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2496 (.out1(_2417), .in1(leafvec82_3629_D), .in2(R12646));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2485 (.out1(_2406), .in1(leafvec82_3629_D), .in2(R12647));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2478 (.out1(_2399), .in1(leafvec82_3629_D), .in2(R12648));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2418 (.out1(_2342), .in1(leafvec88_3637_D), .in2(R12650));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2398 (.out1(_2322), .in1(leafvec88_3637_D), .in2(R12651));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2387 (.out1(_2311), .in1(leafvec88_3637_D), .in2(R12652));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2380 (.out1(_2304), .in1(leafvec88_3637_D), .in2(R12653));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2320 (.out1(_2247), .in1(leafvec94_3645_D), .in2(R12655));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2300 (.out1(_2227), .in1(leafvec94_3645_D), .in2(R12656));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2289 (.out1(_2216), .in1(leafvec94_3645_D), .in2(R12657));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2282 (.out1(_2209), .in1(leafvec94_3645_D), .in2(R12658));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2222 (.out1(_2152), .in1(leafvec100_3653_D), .in2(R12660));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2202 (.out1(_2132), .in1(leafvec100_3653_D), .in2(R12661));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2191 (.out1(_2121), .in1(leafvec100_3653_D), .in2(R12662));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2184 (.out1(_2114), .in1(leafvec100_3653_D), .in2(R12663));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2124 (.out1(_2057), .in1(leafvec106_3661_D), .in2(R12665));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2104 (.out1(_2037), .in1(leafvec106_3661_D), .in2(R12666));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2093 (.out1(_2026), .in1(leafvec106_3661_D), .in2(R12667));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2086 (.out1(_2019), .in1(leafvec106_3661_D), .in2(R12668));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2026 (.out1(_1962), .in1(leafvec112_3669_D), .in2(R12670));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2006 (.out1(_1942), .in1(leafvec112_3669_D), .in2(R12671));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1995 (.out1(_1931), .in1(leafvec112_3669_D), .in2(R12672));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1988 (.out1(_1924), .in1(leafvec112_3669_D), .in2(R12673));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1928 (.out1(_1867), .in1(leafvec118_3677_D), .in2(R12675));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1908 (.out1(_1847), .in1(leafvec118_3677_D), .in2(R12676));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1897 (.out1(_1836), .in1(leafvec118_3677_D), .in2(R12677));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1890 (.out1(_1829), .in1(leafvec118_3677_D), .in2(R12678));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1830 (.out1(_1772), .in1(leafvec124_3684_D), .in2(R12680));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1810 (.out1(_1752), .in1(leafvec124_3684_D), .in2(R12681));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1799 (.out1(_1741), .in1(leafvec124_3684_D), .in2(R12682));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1792 (.out1(_1734), .in1(leafvec124_3684_D), .in2(R12683));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2642 (.out1(_2560), .in1(R12639), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2544 (.out1(_2465), .in1(R12644), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2446 (.out1(_2370), .in1(R12649), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2348 (.out1(_2275), .in1(R12654), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2250 (.out1(_2180), .in1(R12659), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2152 (.out1(_2085), .in1(R12664), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2054 (.out1(_1990), .in1(R12669), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1956 (.out1(_1895), .in1(R12674), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1858 (.out1(_1800), .in1(R12679), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3931 (.out1(R3932), .clock(clock), .in1(R3931));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4187 (.out1(R4188), .clock(clock), .in1(R4187));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4442 (.out1(R4443), .clock(clock), .in1(R4442));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4687 (.out1(R4688), .clock(clock), .in1(R4687));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4927 (.out1(R4928), .clock(clock), .in1(R4927));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5214 (.out1(R5215), .clock(clock), .in1(R5214));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5446 (.out1(R5447), .clock(clock), .in1(R5446));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5673 (.out1(R5674), .clock(clock), .in1(R5673));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5947 (.out1(R5948), .clock(clock), .in1(R5947));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6165 (.out1(R6166), .clock(clock), .in1(R6165));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6378 (.out1(R6379), .clock(clock), .in1(R6378));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6639 (.out1(R6640), .clock(clock), .in1(R6639));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6844 (.out1(R6845), .clock(clock), .in1(R6844));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7044 (.out1(R7045), .clock(clock), .in1(R7044));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7291 (.out1(R7292), .clock(clock), .in1(R7291));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7483 (.out1(R7484), .clock(clock), .in1(R7483));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7670 (.out1(R7671), .clock(clock), .in1(R7670));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7904 (.out1(R7905), .clock(clock), .in1(R7904));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8083 (.out1(R8084), .clock(clock), .in1(R8083));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8257 (.out1(R8258), .clock(clock), .in1(R8257));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8478 (.out1(R8479), .clock(clock), .in1(R8478));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8644 (.out1(R8645), .clock(clock), .in1(R8644));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8805 (.out1(R8806), .clock(clock), .in1(R8805));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9013 (.out1(R9014), .clock(clock), .in1(R9013));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9166 (.out1(R9167), .clock(clock), .in1(R9166));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9314 (.out1(R9315), .clock(clock), .in1(R9314));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9509 (.out1(R9510), .clock(clock), .in1(R9509));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9649 (.out1(R9650), .clock(clock), .in1(R9649));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9784 (.out1(R9785), .clock(clock), .in1(R9784));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9966 (.out1(R9967), .clock(clock), .in1(R9966));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10093 (.out1(R10094), .clock(clock), .in1(R10093));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10215 (.out1(R10216), .clock(clock), .in1(R10215));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10384 (.out1(R10385), .clock(clock), .in1(R10384));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10497 (.out1(R10498), .clock(clock), .in1(R10497));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10605 (.out1(R10606), .clock(clock), .in1(R10605));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10761 (.out1(R10762), .clock(clock), .in1(R10761));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10861 (.out1(R10862), .clock(clock), .in1(R10861));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10956 (.out1(R10957), .clock(clock), .in1(R10956));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11098 (.out1(R11099), .clock(clock), .in1(R11098));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11185 (.out1(R11186), .clock(clock), .in1(R11185));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11267 (.out1(R11268), .clock(clock), .in1(R11267));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11396 (.out1(R11397), .clock(clock), .in1(R11396));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11470 (.out1(R11471), .clock(clock), .in1(R11470));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11539 (.out1(R11540), .clock(clock), .in1(R11539));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11655 (.out1(R11656), .clock(clock), .in1(R11655));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11716 (.out1(R11717), .clock(clock), .in1(R11716));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11772 (.out1(R11773), .clock(clock), .in1(R11772));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11875 (.out1(R11876), .clock(clock), .in1(R11875));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11923 (.out1(R11924), .clock(clock), .in1(R11923));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11966 (.out1(R11967), .clock(clock), .in1(R11966));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12056 (.out1(R12057), .clock(clock), .in1(R12056));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12091 (.out1(R12092), .clock(clock), .in1(R12091));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12121 (.out1(R12122), .clock(clock), .in1(R12121));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12198 (.out1(R12199), .clock(clock), .in1(R12198));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12220 (.out1(R12221), .clock(clock), .in1(R12220));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12237 (.out1(R12238), .clock(clock), .in1(R12237));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12301 (.out1(R12302), .clock(clock), .in1(R12301));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12363 (.out1(R12364), .clock(clock), .in1(R12363));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12377 (.out1(R12378), .clock(clock), .in1(R12377));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12388 (.out1(R12389), .clock(clock), .in1(R12388));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12399 (.out1(R12400), .clock(clock), .in1(R12399));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12410 (.out1(R12411), .clock(clock), .in1(R12410));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12421 (.out1(R12422), .clock(clock), .in1(R12421));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12432 (.out1(R12433), .clock(clock), .in1(R12432));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12443 (.out1(R12444), .clock(clock), .in1(R12443));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12454 (.out1(R12455), .clock(clock), .in1(R12454));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12465 (.out1(R12466), .clock(clock), .in1(R12465));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12519 (.out1(R12520), .clock(clock), .in1(R12519));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12530 (.out1(R12531), .clock(clock), .in1(R12530));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12541 (.out1(R12542), .clock(clock), .in1(R12541));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12552 (.out1(R12553), .clock(clock), .in1(R12552));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12563 (.out1(R12564), .clock(clock), .in1(R12563));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12574 (.out1(R12575), .clock(clock), .in1(R12574));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12585 (.out1(R12586), .clock(clock), .in1(R12585));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12596 (.out1(R12597), .clock(clock), .in1(R12596));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12721 (.out1(R12722), .clock(clock), .in1(_2558));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12722 (.out1(R12723), .clock(clock), .in1(_2551));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12723 (.out1(R12724), .clock(clock), .in1(_2540));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12724 (.out1(R12725), .clock(clock), .in1(_2520));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12725 (.out1(R12726), .clock(clock), .in1(_2463));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12726 (.out1(R12727), .clock(clock), .in1(_2456));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12727 (.out1(R12728), .clock(clock), .in1(_2445));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12728 (.out1(R12729), .clock(clock), .in1(_2425));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12729 (.out1(R12730), .clock(clock), .in1(_2368));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12730 (.out1(R12731), .clock(clock), .in1(_2361));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12731 (.out1(R12732), .clock(clock), .in1(_2350));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12732 (.out1(R12733), .clock(clock), .in1(_2330));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12733 (.out1(R12734), .clock(clock), .in1(_2273));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12734 (.out1(R12735), .clock(clock), .in1(_2266));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12735 (.out1(R12736), .clock(clock), .in1(_2255));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12736 (.out1(R12737), .clock(clock), .in1(_2235));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12737 (.out1(R12738), .clock(clock), .in1(_2178));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12738 (.out1(R12739), .clock(clock), .in1(_2171));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12739 (.out1(R12740), .clock(clock), .in1(_2160));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12740 (.out1(R12741), .clock(clock), .in1(_2140));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12741 (.out1(R12742), .clock(clock), .in1(_2083));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12742 (.out1(R12743), .clock(clock), .in1(_2076));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12743 (.out1(R12744), .clock(clock), .in1(_2065));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12744 (.out1(R12745), .clock(clock), .in1(_2045));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12745 (.out1(R12746), .clock(clock), .in1(_1988));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12746 (.out1(R12747), .clock(clock), .in1(_1981));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12747 (.out1(R12748), .clock(clock), .in1(_1970));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12748 (.out1(R12749), .clock(clock), .in1(_1950));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12749 (.out1(R12750), .clock(clock), .in1(_1893));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12750 (.out1(R12751), .clock(clock), .in1(_1886));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12751 (.out1(R12752), .clock(clock), .in1(_1875));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12752 (.out1(R12753), .clock(clock), .in1(_1855));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12753 (.out1(R12754), .clock(clock), .in1(_1798));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12754 (.out1(R12755), .clock(clock), .in1(_1791));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12755 (.out1(R12756), .clock(clock), .in1(_1780));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12756 (.out1(R12757), .clock(clock), .in1(_1760));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12757 (.out1(R12758), .clock(clock), .in1(ifout3549));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12768 (.out1(R12769), .clock(clock), .in1(ifout3451));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12779 (.out1(R12780), .clock(clock), .in1(_3506));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12780 (.out1(R12781), .clock(clock), .in1(_3499));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12781 (.out1(R12782), .clock(clock), .in1(_3488));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12782 (.out1(R12783), .clock(clock), .in1(_3468));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12783 (.out1(R12784), .clock(clock), .in1(_3411));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12784 (.out1(R12785), .clock(clock), .in1(_3404));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12785 (.out1(R12786), .clock(clock), .in1(_3393));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12786 (.out1(R12787), .clock(clock), .in1(_3373));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12787 (.out1(R12788), .clock(clock), .in1(_3319));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12788 (.out1(R12789), .clock(clock), .in1(_3291));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12789 (.out1(R12790), .clock(clock), .in1(_3271));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12790 (.out1(R12791), .clock(clock), .in1(_3260));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12791 (.out1(R12792), .clock(clock), .in1(_3253));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12792 (.out1(R12793), .clock(clock), .in1(_3224));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12793 (.out1(R12794), .clock(clock), .in1(_3196));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12794 (.out1(R12795), .clock(clock), .in1(_3176));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12795 (.out1(R12796), .clock(clock), .in1(_3165));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12796 (.out1(R12797), .clock(clock), .in1(_3158));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12797 (.out1(R12798), .clock(clock), .in1(_3129));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12798 (.out1(R12799), .clock(clock), .in1(_3101));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12799 (.out1(R12800), .clock(clock), .in1(_3081));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12800 (.out1(R12801), .clock(clock), .in1(_3070));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12801 (.out1(R12802), .clock(clock), .in1(_3063));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12802 (.out1(R12803), .clock(clock), .in1(_3034));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12803 (.out1(R12804), .clock(clock), .in1(_3006));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12804 (.out1(R12805), .clock(clock), .in1(_2986));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12805 (.out1(R12806), .clock(clock), .in1(_2975));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12806 (.out1(R12807), .clock(clock), .in1(_2968));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12807 (.out1(R12808), .clock(clock), .in1(_2939));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12808 (.out1(R12809), .clock(clock), .in1(_2911));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12809 (.out1(R12810), .clock(clock), .in1(_2891));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12810 (.out1(R12811), .clock(clock), .in1(_2880));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12811 (.out1(R12812), .clock(clock), .in1(_2873));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12812 (.out1(R12813), .clock(clock), .in1(_2844));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12813 (.out1(R12814), .clock(clock), .in1(_2816));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12814 (.out1(R12815), .clock(clock), .in1(_2796));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12815 (.out1(R12816), .clock(clock), .in1(_2785));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12816 (.out1(R12817), .clock(clock), .in1(_2778));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12817 (.out1(R12818), .clock(clock), .in1(_2749));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12818 (.out1(R12819), .clock(clock), .in1(_2721));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12819 (.out1(R12820), .clock(clock), .in1(_2701));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12820 (.out1(R12821), .clock(clock), .in1(_2690));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12821 (.out1(R12822), .clock(clock), .in1(_2683));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12822 (.out1(R12823), .clock(clock), .in1(_2654));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12823 (.out1(R12824), .clock(clock), .in1(_2626));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12824 (.out1(R12825), .clock(clock), .in1(_2606));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12825 (.out1(R12826), .clock(clock), .in1(_2595));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12826 (.out1(R12827), .clock(clock), .in1(_2588));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12827 (.out1(R12828), .clock(clock), .in1(_2552));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12828 (.out1(R12829), .clock(clock), .in1(_2541));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12829 (.out1(R12830), .clock(clock), .in1(_2534));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12830 (.out1(R12831), .clock(clock), .in1(_2521));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12831 (.out1(R12832), .clock(clock), .in1(_2514));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12832 (.out1(R12833), .clock(clock), .in1(_2503));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12833 (.out1(R12834), .clock(clock), .in1(_2457));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12834 (.out1(R12835), .clock(clock), .in1(_2446));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12835 (.out1(R12836), .clock(clock), .in1(_2439));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12836 (.out1(R12837), .clock(clock), .in1(_2426));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12837 (.out1(R12838), .clock(clock), .in1(_2419));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12838 (.out1(R12839), .clock(clock), .in1(_2408));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12839 (.out1(R12840), .clock(clock), .in1(_2362));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12840 (.out1(R12841), .clock(clock), .in1(_2351));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12841 (.out1(R12842), .clock(clock), .in1(_2344));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12842 (.out1(R12843), .clock(clock), .in1(_2331));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12843 (.out1(R12844), .clock(clock), .in1(_2324));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12844 (.out1(R12845), .clock(clock), .in1(_2313));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12845 (.out1(R12846), .clock(clock), .in1(_2267));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12846 (.out1(R12847), .clock(clock), .in1(_2256));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12847 (.out1(R12848), .clock(clock), .in1(_2249));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12848 (.out1(R12849), .clock(clock), .in1(_2236));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12849 (.out1(R12850), .clock(clock), .in1(_2229));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12850 (.out1(R12851), .clock(clock), .in1(_2218));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12851 (.out1(R12852), .clock(clock), .in1(_2172));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12852 (.out1(R12853), .clock(clock), .in1(_2161));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12853 (.out1(R12854), .clock(clock), .in1(_2154));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12854 (.out1(R12855), .clock(clock), .in1(_2141));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12855 (.out1(R12856), .clock(clock), .in1(_2134));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12856 (.out1(R12857), .clock(clock), .in1(_2123));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12857 (.out1(R12858), .clock(clock), .in1(_2077));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12858 (.out1(R12859), .clock(clock), .in1(_2066));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12859 (.out1(R12860), .clock(clock), .in1(_2059));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12860 (.out1(R12861), .clock(clock), .in1(_2046));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12861 (.out1(R12862), .clock(clock), .in1(_2039));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12862 (.out1(R12863), .clock(clock), .in1(_2028));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12863 (.out1(R12864), .clock(clock), .in1(_1982));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12864 (.out1(R12865), .clock(clock), .in1(_1971));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12865 (.out1(R12866), .clock(clock), .in1(_1964));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12866 (.out1(R12867), .clock(clock), .in1(_1951));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12867 (.out1(R12868), .clock(clock), .in1(_1944));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12868 (.out1(R12869), .clock(clock), .in1(_1933));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12869 (.out1(R12870), .clock(clock), .in1(_1887));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12870 (.out1(R12871), .clock(clock), .in1(_1876));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12871 (.out1(R12872), .clock(clock), .in1(_1869));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12872 (.out1(R12873), .clock(clock), .in1(_1856));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12873 (.out1(R12874), .clock(clock), .in1(_1849));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12874 (.out1(R12875), .clock(clock), .in1(_1838));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12875 (.out1(R12876), .clock(clock), .in1(_1792));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12876 (.out1(R12877), .clock(clock), .in1(_1781));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12877 (.out1(R12878), .clock(clock), .in1(_1774));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12878 (.out1(R12879), .clock(clock), .in1(_1761));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12879 (.out1(R12880), .clock(clock), .in1(_1754));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12880 (.out1(R12881), .clock(clock), .in1(_1743));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12881 (.out1(R12882), .clock(clock), .in1(_3317));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12882 (.out1(R12883), .clock(clock), .in1(_3310));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12883 (.out1(R12884), .clock(clock), .in1(_3299));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12884 (.out1(R12885), .clock(clock), .in1(_3279));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12885 (.out1(R12886), .clock(clock), .in1(_3222));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12886 (.out1(R12887), .clock(clock), .in1(_3215));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12887 (.out1(R12888), .clock(clock), .in1(_3204));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12888 (.out1(R12889), .clock(clock), .in1(_3184));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12889 (.out1(R12890), .clock(clock), .in1(_3127));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12890 (.out1(R12891), .clock(clock), .in1(_3120));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12891 (.out1(R12892), .clock(clock), .in1(_3109));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12892 (.out1(R12893), .clock(clock), .in1(_3089));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12893 (.out1(R12894), .clock(clock), .in1(_3032));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12894 (.out1(R12895), .clock(clock), .in1(_3025));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12895 (.out1(R12896), .clock(clock), .in1(_3014));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12896 (.out1(R12897), .clock(clock), .in1(_2994));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12897 (.out1(R12898), .clock(clock), .in1(_2937));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12898 (.out1(R12899), .clock(clock), .in1(_2930));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12899 (.out1(R12900), .clock(clock), .in1(_2919));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12900 (.out1(R12901), .clock(clock), .in1(_2899));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12901 (.out1(R12902), .clock(clock), .in1(_2842));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12902 (.out1(R12903), .clock(clock), .in1(_2835));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12903 (.out1(R12904), .clock(clock), .in1(_2824));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12904 (.out1(R12905), .clock(clock), .in1(_2804));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12905 (.out1(R12906), .clock(clock), .in1(_2747));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12906 (.out1(R12907), .clock(clock), .in1(_2740));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12907 (.out1(R12908), .clock(clock), .in1(_2729));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12908 (.out1(R12909), .clock(clock), .in1(_2709));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12909 (.out1(R12910), .clock(clock), .in1(_2652));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12910 (.out1(R12911), .clock(clock), .in1(_2645));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12911 (.out1(R12912), .clock(clock), .in1(_2634));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12912 (.out1(R12913), .clock(clock), .in1(_2614));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12913 (.out1(R12914), .clock(clock), .in1(_2532));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12914 (.out1(R12915), .clock(clock), .in1(_2512));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12915 (.out1(R12916), .clock(clock), .in1(_2501));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12916 (.out1(R12917), .clock(clock), .in1(_2494));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12917 (.out1(R12918), .clock(clock), .in1(_2437));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12918 (.out1(R12919), .clock(clock), .in1(_2417));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12919 (.out1(R12920), .clock(clock), .in1(_2406));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12920 (.out1(R12921), .clock(clock), .in1(_2399));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12921 (.out1(R12922), .clock(clock), .in1(_2342));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12922 (.out1(R12923), .clock(clock), .in1(_2322));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12923 (.out1(R12924), .clock(clock), .in1(_2311));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12924 (.out1(R12925), .clock(clock), .in1(_2304));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12925 (.out1(R12926), .clock(clock), .in1(_2247));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12926 (.out1(R12927), .clock(clock), .in1(_2227));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12927 (.out1(R12928), .clock(clock), .in1(_2216));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12928 (.out1(R12929), .clock(clock), .in1(_2209));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12929 (.out1(R12930), .clock(clock), .in1(_2152));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12930 (.out1(R12931), .clock(clock), .in1(_2132));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12931 (.out1(R12932), .clock(clock), .in1(_2121));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12932 (.out1(R12933), .clock(clock), .in1(_2114));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12933 (.out1(R12934), .clock(clock), .in1(_2057));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12934 (.out1(R12935), .clock(clock), .in1(_2037));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12935 (.out1(R12936), .clock(clock), .in1(_2026));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12936 (.out1(R12937), .clock(clock), .in1(_2019));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12937 (.out1(R12938), .clock(clock), .in1(_1962));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12938 (.out1(R12939), .clock(clock), .in1(_1942));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12939 (.out1(R12940), .clock(clock), .in1(_1931));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12940 (.out1(R12941), .clock(clock), .in1(_1924));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12941 (.out1(R12942), .clock(clock), .in1(_1867));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12942 (.out1(R12943), .clock(clock), .in1(_1847));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12943 (.out1(R12944), .clock(clock), .in1(_1836));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12944 (.out1(R12945), .clock(clock), .in1(_1829));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12945 (.out1(R12946), .clock(clock), .in1(_1772));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12946 (.out1(R12947), .clock(clock), .in1(_1752));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12947 (.out1(R12948), .clock(clock), .in1(_1741));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12948 (.out1(R12949), .clock(clock), .in1(_1734));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12949 (.out1(R12950), .clock(clock), .in1(_2560));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12950 (.out1(R12951), .clock(clock), .in1(_2465));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12951 (.out1(R12952), .clock(clock), .in1(_2370));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12952 (.out1(R12953), .clock(clock), .in1(_2275));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12953 (.out1(R12954), .clock(clock), .in1(_2180));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12954 (.out1(R12955), .clock(clock), .in1(_2085));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12955 (.out1(R12956), .clock(clock), .in1(_1990));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12956 (.out1(R12957), .clock(clock), .in1(_1895));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12957 (.out1(R12958), .clock(clock), .in1(_1800));
  SRAM op3424 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3318),.ADR(R12882));
  SRAM op3417 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3311),.ADR(R12883));
  SRAM op3406 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3300),.ADR(R12884));
  SRAM op3386 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3280),.ADR(R12885));
  SRAM op3326 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3223),.ADR(R12886));
  SRAM op3319 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3216),.ADR(R12887));
  SRAM op3308 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3205),.ADR(R12888));
  SRAM op3288 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3185),.ADR(R12889));
  SRAM op3228 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3128),.ADR(R12890));
  SRAM op3221 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3121),.ADR(R12891));
  SRAM op3210 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3110),.ADR(R12892));
  SRAM op3190 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3090),.ADR(R12893));
  SRAM op3130 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3033),.ADR(R12894));
  SRAM op3123 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3026),.ADR(R12895));
  SRAM op3112 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3015),.ADR(R12896));
  SRAM op3092 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2995),.ADR(R12897));
  SRAM op3032 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2938),.ADR(R12898));
  SRAM op3025 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2931),.ADR(R12899));
  SRAM op3014 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2920),.ADR(R12900));
  SRAM op2994 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2900),.ADR(R12901));
  SRAM op2934 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2843),.ADR(R12902));
  SRAM op2927 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2836),.ADR(R12903));
  SRAM op2916 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2825),.ADR(R12904));
  SRAM op2896 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2805),.ADR(R12905));
  SRAM op2836 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2748),.ADR(R12906));
  SRAM op2829 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2741),.ADR(R12907));
  SRAM op2818 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2730),.ADR(R12908));
  SRAM op2798 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2710),.ADR(R12909));
  SRAM op2738 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2653),.ADR(R12910));
  SRAM op2731 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2646),.ADR(R12911));
  SRAM op2720 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2635),.ADR(R12912));
  SRAM op2700 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2615),.ADR(R12913));
  SRAM op2615 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2533),.ADR(R12914));
  SRAM op2595 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2513),.ADR(R12915));
  SRAM op2584 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2502),.ADR(R12916));
  SRAM op2577 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2495),.ADR(R12917));
  SRAM op2517 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2438),.ADR(R12918));
  SRAM op2497 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2418),.ADR(R12919));
  SRAM op2486 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2407),.ADR(R12920));
  SRAM op2479 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2400),.ADR(R12921));
  SRAM op2419 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2343),.ADR(R12922));
  SRAM op2399 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2323),.ADR(R12923));
  SRAM op2388 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2312),.ADR(R12924));
  SRAM op2381 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2305),.ADR(R12925));
  SRAM op2321 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2248),.ADR(R12926));
  SRAM op2301 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2228),.ADR(R12927));
  SRAM op2290 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2217),.ADR(R12928));
  SRAM op2283 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2210),.ADR(R12929));
  SRAM op2223 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2153),.ADR(R12930));
  SRAM op2203 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2133),.ADR(R12931));
  SRAM op2192 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2122),.ADR(R12932));
  SRAM op2185 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2115),.ADR(R12933));
  SRAM op2125 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2058),.ADR(R12934));
  SRAM op2105 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2038),.ADR(R12935));
  SRAM op2094 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2027),.ADR(R12936));
  SRAM op2087 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2020),.ADR(R12937));
  SRAM op2027 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1963),.ADR(R12938));
  SRAM op2007 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1943),.ADR(R12939));
  SRAM op1996 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1932),.ADR(R12940));
  SRAM op1989 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1925),.ADR(R12941));
  SRAM op1929 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1868),.ADR(R12942));
  SRAM op1909 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1848),.ADR(R12943));
  SRAM op1898 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1837),.ADR(R12944));
  SRAM op1891 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1830),.ADR(R12945));
  SRAM op1831 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1773),.ADR(R12946));
  SRAM op1811 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1753),.ADR(R12947));
  SRAM op1800 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1742),.ADR(R12948));
  SRAM op1793 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1735),.ADR(R12949));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3592 (.out1(_3480), .in1(R4443));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3572 (.out1(_3460), .in1(R4443));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3561 (.out1(_3449), .in1(R4443));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3554 (.out1(_3442), .in1(R4443));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3494 (.out1(_3385), .in1(R5215));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3474 (.out1(_3365), .in1(R5215));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3463 (.out1(_3354), .in1(R5215));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3456 (.out1(_3347), .in1(R5215));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2643 (.out1(_2561), .in1(R12722), .in2(R12950));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2545 (.out1(_2466), .in1(R12726), .in2(R12951));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2447 (.out1(_2371), .in1(R12730), .in2(R12952));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2349 (.out1(_2276), .in1(R12734), .in2(R12953));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2251 (.out1(_2181), .in1(R12738), .in2(R12954));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2153 (.out1(_2086), .in1(R12742), .in2(R12955));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2055 (.out1(_1991), .in1(R12746), .in2(R12956));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1957 (.out1(_1896), .in1(R12750), .in2(R12957));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1859 (.out1(_1801), .in1(R12754), .in2(R12958));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2644 (.out1(_2562), .in1(_2561), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2635 (.out1(_2553), .in1(R12828), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2624 (.out1(_2542), .in1(R12829), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2604 (.out1(_2522), .in1(R12831), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2546 (.out1(_2467), .in1(_2466), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2537 (.out1(_2458), .in1(R12834), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2526 (.out1(_2447), .in1(R12835), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2506 (.out1(_2427), .in1(R12837), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2448 (.out1(_2372), .in1(_2371), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2439 (.out1(_2363), .in1(R12840), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2428 (.out1(_2352), .in1(R12841), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2408 (.out1(_2332), .in1(R12843), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2350 (.out1(_2277), .in1(_2276), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2341 (.out1(_2268), .in1(R12846), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2330 (.out1(_2257), .in1(R12847), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2310 (.out1(_2237), .in1(R12849), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2252 (.out1(_2182), .in1(_2181), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2243 (.out1(_2173), .in1(R12852), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2232 (.out1(_2162), .in1(R12853), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2212 (.out1(_2142), .in1(R12855), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2154 (.out1(_2087), .in1(_2086), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2145 (.out1(_2078), .in1(R12858), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2134 (.out1(_2067), .in1(R12859), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2114 (.out1(_2047), .in1(R12861), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2056 (.out1(_1992), .in1(_1991), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2047 (.out1(_1983), .in1(R12864), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2036 (.out1(_1972), .in1(R12865), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2016 (.out1(_1952), .in1(R12867), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1958 (.out1(_1897), .in1(_1896), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1949 (.out1(_1888), .in1(R12870), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1938 (.out1(_1877), .in1(R12871), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1918 (.out1(_1857), .in1(R12873), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1860 (.out1(_1802), .in1(_1801), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1851 (.out1(_1793), .in1(R12876), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1840 (.out1(_1782), .in1(R12877), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1820 (.out1(_1762), .in1(R12879), .in2(64 'd 18446744073709551615));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3621 (.out1(_3509), .in1(2 'd 2), .in2(R4688));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3593 (.out1(_3481), .in1(_3480), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3573 (.out1(_3461), .in1(_3460), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3562 (.out1(_3450), .in1(_3449), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3555 (.out1(_3443), .in1(_3442), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3523 (.out1(_3414), .in1(2 'd 2), .in2(R5447));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3495 (.out1(_3386), .in1(_3385), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3475 (.out1(_3366), .in1(_3365), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3464 (.out1(_3355), .in1(_3354), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3457 (.out1(_3348), .in1(_3347), .in2(2 'd 3));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3418 (.out1(_3312), .in1(2 'd 2), .in2(R6166));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3407 (.out1(_3301), .in1(2 'd 2), .in2(R6166));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3400 (.out1(_3294), .in1(2 'd 2), .in2(R6166));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3387 (.out1(_3281), .in1(2 'd 2), .in2(R6166));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3380 (.out1(_3274), .in1(2 'd 2), .in2(R6166));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3369 (.out1(_3263), .in1(2 'd 2), .in2(R6166));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3320 (.out1(_3217), .in1(2 'd 2), .in2(R6845));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3309 (.out1(_3206), .in1(2 'd 2), .in2(R6845));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3302 (.out1(_3199), .in1(2 'd 2), .in2(R6845));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3289 (.out1(_3186), .in1(2 'd 2), .in2(R6845));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3282 (.out1(_3179), .in1(2 'd 2), .in2(R6845));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3271 (.out1(_3168), .in1(2 'd 2), .in2(R6845));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3222 (.out1(_3122), .in1(2 'd 2), .in2(R7484));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3211 (.out1(_3111), .in1(2 'd 2), .in2(R7484));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3204 (.out1(_3104), .in1(2 'd 2), .in2(R7484));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3191 (.out1(_3091), .in1(2 'd 2), .in2(R7484));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3184 (.out1(_3084), .in1(2 'd 2), .in2(R7484));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3173 (.out1(_3073), .in1(2 'd 2), .in2(R7484));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3124 (.out1(_3027), .in1(2 'd 2), .in2(R8084));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3113 (.out1(_3016), .in1(2 'd 2), .in2(R8084));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3106 (.out1(_3009), .in1(2 'd 2), .in2(R8084));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3093 (.out1(_2996), .in1(2 'd 2), .in2(R8084));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3086 (.out1(_2989), .in1(2 'd 2), .in2(R8084));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3075 (.out1(_2978), .in1(2 'd 2), .in2(R8084));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3026 (.out1(_2932), .in1(2 'd 2), .in2(R8645));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3015 (.out1(_2921), .in1(2 'd 2), .in2(R8645));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3008 (.out1(_2914), .in1(2 'd 2), .in2(R8645));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2995 (.out1(_2901), .in1(2 'd 2), .in2(R8645));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2988 (.out1(_2894), .in1(2 'd 2), .in2(R8645));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2977 (.out1(_2883), .in1(2 'd 2), .in2(R8645));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2928 (.out1(_2837), .in1(2 'd 2), .in2(R9167));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2917 (.out1(_2826), .in1(2 'd 2), .in2(R9167));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2910 (.out1(_2819), .in1(2 'd 2), .in2(R9167));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2897 (.out1(_2806), .in1(2 'd 2), .in2(R9167));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2890 (.out1(_2799), .in1(2 'd 2), .in2(R9167));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2879 (.out1(_2788), .in1(2 'd 2), .in2(R9167));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2830 (.out1(_2742), .in1(2 'd 2), .in2(R9650));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2819 (.out1(_2731), .in1(2 'd 2), .in2(R9650));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2812 (.out1(_2724), .in1(2 'd 2), .in2(R9650));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2799 (.out1(_2711), .in1(2 'd 2), .in2(R9650));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2792 (.out1(_2704), .in1(2 'd 2), .in2(R9650));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2781 (.out1(_2693), .in1(2 'd 2), .in2(R9650));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2732 (.out1(_2647), .in1(2 'd 2), .in2(R10094));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2721 (.out1(_2636), .in1(2 'd 2), .in2(R10094));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2714 (.out1(_2629), .in1(2 'd 2), .in2(R10094));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2701 (.out1(_2616), .in1(2 'd 2), .in2(R10094));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2694 (.out1(_2609), .in1(2 'd 2), .in2(R10094));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2683 (.out1(_2598), .in1(2 'd 2), .in2(R10094));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2578 (.out1(_2496), .in1(2 'd 2), .in2(R10498));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2480 (.out1(_2401), .in1(2 'd 2), .in2(R10862));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2382 (.out1(_2306), .in1(2 'd 2), .in2(R11186));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2284 (.out1(_2211), .in1(2 'd 2), .in2(R11471));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2186 (.out1(_2116), .in1(2 'd 2), .in2(R11717));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2088 (.out1(_2021), .in1(2 'd 2), .in2(R11924));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1990 (.out1(_1926), .in1(2 'd 2), .in2(R12092));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1892 (.out1(_1831), .in1(2 'd 2), .in2(R12221));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op1794 (.out1(_1736), .in1(2 'd 2), .in2(R12364));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3619 (.out1(_3507), .in1(leafvec16_3539_D), .in2(R12780));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3612 (.out1(_3500), .in1(leafvec16_3539_D), .in2(R12781));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3601 (.out1(_3489), .in1(leafvec16_3539_D), .in2(R12782));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3581 (.out1(_3469), .in1(leafvec16_3539_D), .in2(R12783));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3521 (.out1(_3412), .in1(leafvec22_3548_D), .in2(R12784));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3514 (.out1(_3405), .in1(leafvec22_3548_D), .in2(R12785));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3503 (.out1(_3394), .in1(leafvec22_3548_D), .in2(R12786));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3483 (.out1(_3374), .in1(leafvec22_3548_D), .in2(R12787));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3398 (.out1(_3292), .in1(leafvec28_3556_D), .in2(R12789));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3378 (.out1(_3272), .in1(leafvec28_3556_D), .in2(R12790));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3367 (.out1(_3261), .in1(leafvec28_3556_D), .in2(R12791));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3360 (.out1(_3254), .in1(leafvec28_3556_D), .in2(R12792));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3300 (.out1(_3197), .in1(leafvec34_3564_D), .in2(R12794));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3280 (.out1(_3177), .in1(leafvec34_3564_D), .in2(R12795));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3269 (.out1(_3166), .in1(leafvec34_3564_D), .in2(R12796));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3262 (.out1(_3159), .in1(leafvec34_3564_D), .in2(R12797));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3202 (.out1(_3102), .in1(leafvec40_3572_D), .in2(R12799));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3182 (.out1(_3082), .in1(leafvec40_3572_D), .in2(R12800));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3171 (.out1(_3071), .in1(leafvec40_3572_D), .in2(R12801));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3164 (.out1(_3064), .in1(leafvec40_3572_D), .in2(R12802));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3104 (.out1(_3007), .in1(leafvec46_3580_D), .in2(R12804));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3084 (.out1(_2987), .in1(leafvec46_3580_D), .in2(R12805));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3073 (.out1(_2976), .in1(leafvec46_3580_D), .in2(R12806));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3066 (.out1(_2969), .in1(leafvec46_3580_D), .in2(R12807));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3006 (.out1(_2912), .in1(leafvec52_3588_D), .in2(R12809));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2986 (.out1(_2892), .in1(leafvec52_3588_D), .in2(R12810));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2975 (.out1(_2881), .in1(leafvec52_3588_D), .in2(R12811));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2968 (.out1(_2874), .in1(leafvec52_3588_D), .in2(R12812));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2908 (.out1(_2817), .in1(leafvec58_3596_D), .in2(R12814));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2888 (.out1(_2797), .in1(leafvec58_3596_D), .in2(R12815));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2877 (.out1(_2786), .in1(leafvec58_3596_D), .in2(R12816));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2870 (.out1(_2779), .in1(leafvec58_3596_D), .in2(R12817));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2810 (.out1(_2722), .in1(leafvec64_3605_D), .in2(R12819));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2790 (.out1(_2702), .in1(leafvec64_3605_D), .in2(R12820));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2779 (.out1(_2691), .in1(leafvec64_3605_D), .in2(R12821));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2772 (.out1(_2684), .in1(leafvec64_3605_D), .in2(R12822));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2712 (.out1(_2627), .in1(leafvec70_3613_D), .in2(R12824));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2692 (.out1(_2607), .in1(leafvec70_3613_D), .in2(R12825));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2681 (.out1(_2596), .in1(leafvec70_3613_D), .in2(R12826));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2674 (.out1(_2589), .in1(leafvec70_3613_D), .in2(R12827));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2645 (.out1(_2563), .in1(_2562), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2636 (.out1(_2554), .in1(R12723), .in2(_2553));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2625 (.out1(_2543), .in1(R12724), .in2(_2542));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2605 (.out1(_2523), .in1(R12725), .in2(_2522));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2547 (.out1(_2468), .in1(_2467), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2538 (.out1(_2459), .in1(R12727), .in2(_2458));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2527 (.out1(_2448), .in1(R12728), .in2(_2447));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2507 (.out1(_2428), .in1(R12729), .in2(_2427));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2449 (.out1(_2373), .in1(_2372), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2440 (.out1(_2364), .in1(R12731), .in2(_2363));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2429 (.out1(_2353), .in1(R12732), .in2(_2352));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2409 (.out1(_2333), .in1(R12733), .in2(_2332));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2351 (.out1(_2278), .in1(_2277), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2342 (.out1(_2269), .in1(R12735), .in2(_2268));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2331 (.out1(_2258), .in1(R12736), .in2(_2257));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2311 (.out1(_2238), .in1(R12737), .in2(_2237));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2253 (.out1(_2183), .in1(_2182), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2244 (.out1(_2174), .in1(R12739), .in2(_2173));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2233 (.out1(_2163), .in1(R12740), .in2(_2162));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2213 (.out1(_2143), .in1(R12741), .in2(_2142));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2155 (.out1(_2088), .in1(_2087), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2146 (.out1(_2079), .in1(R12743), .in2(_2078));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2135 (.out1(_2068), .in1(R12744), .in2(_2067));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2115 (.out1(_2048), .in1(R12745), .in2(_2047));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2057 (.out1(_1993), .in1(_1992), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2048 (.out1(_1984), .in1(R12747), .in2(_1983));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2037 (.out1(_1973), .in1(R12748), .in2(_1972));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2017 (.out1(_1953), .in1(R12749), .in2(_1952));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1959 (.out1(_1898), .in1(_1897), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1950 (.out1(_1889), .in1(R12751), .in2(_1888));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1939 (.out1(_1878), .in1(R12752), .in2(_1877));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1919 (.out1(_1858), .in1(R12753), .in2(_1857));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1861 (.out1(_1803), .in1(_1802), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1852 (.out1(_1794), .in1(R12755), .in2(_1793));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1841 (.out1(_1783), .in1(R12756), .in2(_1782));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1821 (.out1(_1763), .in1(R12757), .in2(_1762));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3426 (.out1(_3320), .in1(R12788), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3328 (.out1(_3225), .in1(R12793), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3230 (.out1(_3130), .in1(R12798), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3132 (.out1(_3035), .in1(R12803), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3034 (.out1(_2940), .in1(R12808), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2936 (.out1(_2845), .in1(R12813), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2838 (.out1(_2750), .in1(R12818), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2740 (.out1(_2655), .in1(R12823), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2646 (.out1(_2564), .in1(_2554), .in2(_2563));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2626 (.out1(_2544), .in1(_2543), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2617 (.out1(_2535), .in1(R12830), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2606 (.out1(_2524), .in1(_2523), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2597 (.out1(_2515), .in1(R12832), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2586 (.out1(_2504), .in1(R12833), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2548 (.out1(_2469), .in1(_2459), .in2(_2468));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2528 (.out1(_2449), .in1(_2448), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2519 (.out1(_2440), .in1(R12836), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2508 (.out1(_2429), .in1(_2428), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2499 (.out1(_2420), .in1(R12838), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2488 (.out1(_2409), .in1(R12839), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2450 (.out1(_2374), .in1(_2364), .in2(_2373));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2430 (.out1(_2354), .in1(_2353), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2421 (.out1(_2345), .in1(R12842), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2410 (.out1(_2334), .in1(_2333), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2401 (.out1(_2325), .in1(R12844), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2390 (.out1(_2314), .in1(R12845), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2352 (.out1(_2279), .in1(_2269), .in2(_2278));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2332 (.out1(_2259), .in1(_2258), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2323 (.out1(_2250), .in1(R12848), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2312 (.out1(_2239), .in1(_2238), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2303 (.out1(_2230), .in1(R12850), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2292 (.out1(_2219), .in1(R12851), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2254 (.out1(_2184), .in1(_2174), .in2(_2183));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2234 (.out1(_2164), .in1(_2163), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2225 (.out1(_2155), .in1(R12854), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2214 (.out1(_2144), .in1(_2143), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2205 (.out1(_2135), .in1(R12856), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2194 (.out1(_2124), .in1(R12857), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2156 (.out1(_2089), .in1(_2079), .in2(_2088));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2136 (.out1(_2069), .in1(_2068), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2127 (.out1(_2060), .in1(R12860), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2116 (.out1(_2049), .in1(_2048), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2107 (.out1(_2040), .in1(R12862), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2096 (.out1(_2029), .in1(R12863), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2058 (.out1(_1994), .in1(_1984), .in2(_1993));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2038 (.out1(_1974), .in1(_1973), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2029 (.out1(_1965), .in1(R12866), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2018 (.out1(_1954), .in1(_1953), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2009 (.out1(_1945), .in1(R12868), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1998 (.out1(_1934), .in1(R12869), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1960 (.out1(_1899), .in1(_1889), .in2(_1898));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1940 (.out1(_1879), .in1(_1878), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1931 (.out1(_1870), .in1(R12872), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1920 (.out1(_1859), .in1(_1858), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1911 (.out1(_1850), .in1(R12874), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1900 (.out1(_1839), .in1(R12875), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1862 (.out1(_1804), .in1(_1794), .in2(_1803));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1842 (.out1(_1784), .in1(_1783), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1833 (.out1(_1775), .in1(R12878), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1822 (.out1(_1764), .in1(_1763), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1813 (.out1(_1755), .in1(R12880), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1802 (.out1(_1744), .in1(R12881), .in2(64 'd 18446744073709551615));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3932 (.out1(R3933), .clock(clock), .in1(R3932));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4188 (.out1(R4189), .clock(clock), .in1(R4188));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4443 (.out1(R4444), .clock(clock), .in1(R4443));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4688 (.out1(R4689), .clock(clock), .in1(R4688));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4928 (.out1(R4929), .clock(clock), .in1(R4928));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5215 (.out1(R5216), .clock(clock), .in1(R5215));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5447 (.out1(R5448), .clock(clock), .in1(R5447));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5674 (.out1(R5675), .clock(clock), .in1(R5674));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5948 (.out1(R5949), .clock(clock), .in1(R5948));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6166 (.out1(R6167), .clock(clock), .in1(R6166));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6379 (.out1(R6380), .clock(clock), .in1(R6379));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6640 (.out1(R6641), .clock(clock), .in1(R6640));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6845 (.out1(R6846), .clock(clock), .in1(R6845));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7045 (.out1(R7046), .clock(clock), .in1(R7045));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7292 (.out1(R7293), .clock(clock), .in1(R7292));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7484 (.out1(R7485), .clock(clock), .in1(R7484));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7671 (.out1(R7672), .clock(clock), .in1(R7671));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7905 (.out1(R7906), .clock(clock), .in1(R7905));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8084 (.out1(R8085), .clock(clock), .in1(R8084));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8258 (.out1(R8259), .clock(clock), .in1(R8258));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8479 (.out1(R8480), .clock(clock), .in1(R8479));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8645 (.out1(R8646), .clock(clock), .in1(R8645));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8806 (.out1(R8807), .clock(clock), .in1(R8806));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9014 (.out1(R9015), .clock(clock), .in1(R9014));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9167 (.out1(R9168), .clock(clock), .in1(R9167));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9315 (.out1(R9316), .clock(clock), .in1(R9315));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9510 (.out1(R9511), .clock(clock), .in1(R9510));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9650 (.out1(R9651), .clock(clock), .in1(R9650));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9785 (.out1(R9786), .clock(clock), .in1(R9785));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9967 (.out1(R9968), .clock(clock), .in1(R9967));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10094 (.out1(R10095), .clock(clock), .in1(R10094));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10216 (.out1(R10217), .clock(clock), .in1(R10216));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10385 (.out1(R10386), .clock(clock), .in1(R10385));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10606 (.out1(R10607), .clock(clock), .in1(R10606));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10762 (.out1(R10763), .clock(clock), .in1(R10762));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10957 (.out1(R10958), .clock(clock), .in1(R10957));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11099 (.out1(R11100), .clock(clock), .in1(R11099));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11268 (.out1(R11269), .clock(clock), .in1(R11268));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11397 (.out1(R11398), .clock(clock), .in1(R11397));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11540 (.out1(R11541), .clock(clock), .in1(R11540));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11656 (.out1(R11657), .clock(clock), .in1(R11656));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11773 (.out1(R11774), .clock(clock), .in1(R11773));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11876 (.out1(R11877), .clock(clock), .in1(R11876));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11967 (.out1(R11968), .clock(clock), .in1(R11967));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12057 (.out1(R12058), .clock(clock), .in1(R12057));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12122 (.out1(R12123), .clock(clock), .in1(R12122));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12199 (.out1(R12200), .clock(clock), .in1(R12199));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12238 (.out1(R12239), .clock(clock), .in1(R12238));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12302 (.out1(R12303), .clock(clock), .in1(R12302));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12378 (.out1(R12379), .clock(clock), .in1(R12378));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12389 (.out1(R12390), .clock(clock), .in1(R12389));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12400 (.out1(R12401), .clock(clock), .in1(R12400));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12411 (.out1(R12412), .clock(clock), .in1(R12411));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12422 (.out1(R12423), .clock(clock), .in1(R12422));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12433 (.out1(R12434), .clock(clock), .in1(R12433));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12444 (.out1(R12445), .clock(clock), .in1(R12444));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12455 (.out1(R12456), .clock(clock), .in1(R12455));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12466 (.out1(R12467), .clock(clock), .in1(R12466));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12520 (.out1(R12521), .clock(clock), .in1(R12520));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12531 (.out1(R12532), .clock(clock), .in1(R12531));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12542 (.out1(R12543), .clock(clock), .in1(R12542));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12553 (.out1(R12554), .clock(clock), .in1(R12553));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12564 (.out1(R12565), .clock(clock), .in1(R12564));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12575 (.out1(R12576), .clock(clock), .in1(R12575));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12586 (.out1(R12587), .clock(clock), .in1(R12586));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12597 (.out1(R12598), .clock(clock), .in1(R12597));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12758 (.out1(R12759), .clock(clock), .in1(R12758));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12769 (.out1(R12770), .clock(clock), .in1(R12769));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12958 (.out1(R12959), .clock(clock), .in1(_3318));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12959 (.out1(R12960), .clock(clock), .in1(_3311));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12960 (.out1(R12961), .clock(clock), .in1(_3300));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12961 (.out1(R12962), .clock(clock), .in1(_3280));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12962 (.out1(R12963), .clock(clock), .in1(_3223));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12963 (.out1(R12964), .clock(clock), .in1(_3216));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12964 (.out1(R12965), .clock(clock), .in1(_3205));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12965 (.out1(R12966), .clock(clock), .in1(_3185));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12966 (.out1(R12967), .clock(clock), .in1(_3128));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12967 (.out1(R12968), .clock(clock), .in1(_3121));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12968 (.out1(R12969), .clock(clock), .in1(_3110));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12969 (.out1(R12970), .clock(clock), .in1(_3090));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12970 (.out1(R12971), .clock(clock), .in1(_3033));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12971 (.out1(R12972), .clock(clock), .in1(_3026));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12972 (.out1(R12973), .clock(clock), .in1(_3015));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12973 (.out1(R12974), .clock(clock), .in1(_2995));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12974 (.out1(R12975), .clock(clock), .in1(_2938));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12975 (.out1(R12976), .clock(clock), .in1(_2931));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12976 (.out1(R12977), .clock(clock), .in1(_2920));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12977 (.out1(R12978), .clock(clock), .in1(_2900));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12978 (.out1(R12979), .clock(clock), .in1(_2843));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12979 (.out1(R12980), .clock(clock), .in1(_2836));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12980 (.out1(R12981), .clock(clock), .in1(_2825));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12981 (.out1(R12982), .clock(clock), .in1(_2805));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12982 (.out1(R12983), .clock(clock), .in1(_2748));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12983 (.out1(R12984), .clock(clock), .in1(_2741));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12984 (.out1(R12985), .clock(clock), .in1(_2730));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12985 (.out1(R12986), .clock(clock), .in1(_2710));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12986 (.out1(R12987), .clock(clock), .in1(_2653));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12987 (.out1(R12988), .clock(clock), .in1(_2646));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12988 (.out1(R12989), .clock(clock), .in1(_2635));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12989 (.out1(R12990), .clock(clock), .in1(_2615));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12990 (.out1(R12991), .clock(clock), .in1(_2533));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12991 (.out1(R12992), .clock(clock), .in1(_2513));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12992 (.out1(R12993), .clock(clock), .in1(_2502));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12993 (.out1(R12994), .clock(clock), .in1(_2495));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12994 (.out1(R12995), .clock(clock), .in1(_2438));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12995 (.out1(R12996), .clock(clock), .in1(_2418));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12996 (.out1(R12997), .clock(clock), .in1(_2407));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12997 (.out1(R12998), .clock(clock), .in1(_2400));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12998 (.out1(R12999), .clock(clock), .in1(_2343));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op12999 (.out1(R13000), .clock(clock), .in1(_2323));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13000 (.out1(R13001), .clock(clock), .in1(_2312));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13001 (.out1(R13002), .clock(clock), .in1(_2305));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13002 (.out1(R13003), .clock(clock), .in1(_2248));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13003 (.out1(R13004), .clock(clock), .in1(_2228));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13004 (.out1(R13005), .clock(clock), .in1(_2217));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13005 (.out1(R13006), .clock(clock), .in1(_2210));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13006 (.out1(R13007), .clock(clock), .in1(_2153));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13007 (.out1(R13008), .clock(clock), .in1(_2133));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13008 (.out1(R13009), .clock(clock), .in1(_2122));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13009 (.out1(R13010), .clock(clock), .in1(_2115));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13010 (.out1(R13011), .clock(clock), .in1(_2058));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13011 (.out1(R13012), .clock(clock), .in1(_2038));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13012 (.out1(R13013), .clock(clock), .in1(_2027));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13013 (.out1(R13014), .clock(clock), .in1(_2020));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13014 (.out1(R13015), .clock(clock), .in1(_1963));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13015 (.out1(R13016), .clock(clock), .in1(_1943));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13016 (.out1(R13017), .clock(clock), .in1(_1932));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13017 (.out1(R13018), .clock(clock), .in1(_1925));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13018 (.out1(R13019), .clock(clock), .in1(_1868));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13019 (.out1(R13020), .clock(clock), .in1(_1848));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13020 (.out1(R13021), .clock(clock), .in1(_1837));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13021 (.out1(R13022), .clock(clock), .in1(_1830));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13022 (.out1(R13023), .clock(clock), .in1(_1773));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13023 (.out1(R13024), .clock(clock), .in1(_1753));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13024 (.out1(R13025), .clock(clock), .in1(_1742));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13025 (.out1(R13026), .clock(clock), .in1(_1735));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13026 (.out1(R13027), .clock(clock), .in1(_3509));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13027 (.out1(R13028), .clock(clock), .in1(_3481));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13028 (.out1(R13029), .clock(clock), .in1(_3461));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13029 (.out1(R13030), .clock(clock), .in1(_3450));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13030 (.out1(R13031), .clock(clock), .in1(_3443));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13031 (.out1(R13032), .clock(clock), .in1(_3414));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13032 (.out1(R13033), .clock(clock), .in1(_3386));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13033 (.out1(R13034), .clock(clock), .in1(_3366));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13034 (.out1(R13035), .clock(clock), .in1(_3355));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13035 (.out1(R13036), .clock(clock), .in1(_3348));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13036 (.out1(R13037), .clock(clock), .in1(_3312));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13037 (.out1(R13038), .clock(clock), .in1(_3301));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13038 (.out1(R13039), .clock(clock), .in1(_3294));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13039 (.out1(R13040), .clock(clock), .in1(_3281));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13040 (.out1(R13041), .clock(clock), .in1(_3274));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13041 (.out1(R13042), .clock(clock), .in1(_3263));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13042 (.out1(R13043), .clock(clock), .in1(_3217));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13043 (.out1(R13044), .clock(clock), .in1(_3206));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13044 (.out1(R13045), .clock(clock), .in1(_3199));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13045 (.out1(R13046), .clock(clock), .in1(_3186));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13046 (.out1(R13047), .clock(clock), .in1(_3179));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13047 (.out1(R13048), .clock(clock), .in1(_3168));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13048 (.out1(R13049), .clock(clock), .in1(_3122));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13049 (.out1(R13050), .clock(clock), .in1(_3111));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13050 (.out1(R13051), .clock(clock), .in1(_3104));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13051 (.out1(R13052), .clock(clock), .in1(_3091));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13052 (.out1(R13053), .clock(clock), .in1(_3084));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13053 (.out1(R13054), .clock(clock), .in1(_3073));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13054 (.out1(R13055), .clock(clock), .in1(_3027));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13055 (.out1(R13056), .clock(clock), .in1(_3016));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13056 (.out1(R13057), .clock(clock), .in1(_3009));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13057 (.out1(R13058), .clock(clock), .in1(_2996));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13058 (.out1(R13059), .clock(clock), .in1(_2989));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13059 (.out1(R13060), .clock(clock), .in1(_2978));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13060 (.out1(R13061), .clock(clock), .in1(_2932));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13061 (.out1(R13062), .clock(clock), .in1(_2921));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13062 (.out1(R13063), .clock(clock), .in1(_2914));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13063 (.out1(R13064), .clock(clock), .in1(_2901));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13064 (.out1(R13065), .clock(clock), .in1(_2894));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13065 (.out1(R13066), .clock(clock), .in1(_2883));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13066 (.out1(R13067), .clock(clock), .in1(_2837));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13067 (.out1(R13068), .clock(clock), .in1(_2826));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13068 (.out1(R13069), .clock(clock), .in1(_2819));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13069 (.out1(R13070), .clock(clock), .in1(_2806));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13070 (.out1(R13071), .clock(clock), .in1(_2799));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13071 (.out1(R13072), .clock(clock), .in1(_2788));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13072 (.out1(R13073), .clock(clock), .in1(_2742));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13073 (.out1(R13074), .clock(clock), .in1(_2731));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13074 (.out1(R13075), .clock(clock), .in1(_2724));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13075 (.out1(R13076), .clock(clock), .in1(_2711));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13076 (.out1(R13077), .clock(clock), .in1(_2704));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13077 (.out1(R13078), .clock(clock), .in1(_2693));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13078 (.out1(R13079), .clock(clock), .in1(_2647));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13079 (.out1(R13080), .clock(clock), .in1(_2636));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13080 (.out1(R13081), .clock(clock), .in1(_2629));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13081 (.out1(R13082), .clock(clock), .in1(_2616));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13082 (.out1(R13083), .clock(clock), .in1(_2609));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13083 (.out1(R13084), .clock(clock), .in1(_2598));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13084 (.out1(R13085), .clock(clock), .in1(_2496));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13085 (.out1(R13086), .clock(clock), .in1(_2401));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13086 (.out1(R13087), .clock(clock), .in1(_2306));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13087 (.out1(R13088), .clock(clock), .in1(_2211));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13088 (.out1(R13089), .clock(clock), .in1(_2116));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13089 (.out1(R13090), .clock(clock), .in1(_2021));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13090 (.out1(R13091), .clock(clock), .in1(_1926));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13091 (.out1(R13092), .clock(clock), .in1(_1831));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13092 (.out1(R13093), .clock(clock), .in1(_1736));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13093 (.out1(R13094), .clock(clock), .in1(_3507));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13094 (.out1(R13095), .clock(clock), .in1(_3500));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13095 (.out1(R13096), .clock(clock), .in1(_3489));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13096 (.out1(R13097), .clock(clock), .in1(_3469));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13097 (.out1(R13098), .clock(clock), .in1(_3412));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13098 (.out1(R13099), .clock(clock), .in1(_3405));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13099 (.out1(R13100), .clock(clock), .in1(_3394));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13100 (.out1(R13101), .clock(clock), .in1(_3374));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13101 (.out1(R13102), .clock(clock), .in1(_3292));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13102 (.out1(R13103), .clock(clock), .in1(_3272));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13103 (.out1(R13104), .clock(clock), .in1(_3261));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13104 (.out1(R13105), .clock(clock), .in1(_3254));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13105 (.out1(R13106), .clock(clock), .in1(_3197));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13106 (.out1(R13107), .clock(clock), .in1(_3177));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13107 (.out1(R13108), .clock(clock), .in1(_3166));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13108 (.out1(R13109), .clock(clock), .in1(_3159));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13109 (.out1(R13110), .clock(clock), .in1(_3102));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13110 (.out1(R13111), .clock(clock), .in1(_3082));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13111 (.out1(R13112), .clock(clock), .in1(_3071));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13112 (.out1(R13113), .clock(clock), .in1(_3064));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13113 (.out1(R13114), .clock(clock), .in1(_3007));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13114 (.out1(R13115), .clock(clock), .in1(_2987));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13115 (.out1(R13116), .clock(clock), .in1(_2976));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13116 (.out1(R13117), .clock(clock), .in1(_2969));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13117 (.out1(R13118), .clock(clock), .in1(_2912));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13118 (.out1(R13119), .clock(clock), .in1(_2892));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13119 (.out1(R13120), .clock(clock), .in1(_2881));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13120 (.out1(R13121), .clock(clock), .in1(_2874));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13121 (.out1(R13122), .clock(clock), .in1(_2817));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13122 (.out1(R13123), .clock(clock), .in1(_2797));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13123 (.out1(R13124), .clock(clock), .in1(_2786));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13124 (.out1(R13125), .clock(clock), .in1(_2779));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13125 (.out1(R13126), .clock(clock), .in1(_2722));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13126 (.out1(R13127), .clock(clock), .in1(_2702));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13127 (.out1(R13128), .clock(clock), .in1(_2691));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13128 (.out1(R13129), .clock(clock), .in1(_2684));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13129 (.out1(R13130), .clock(clock), .in1(_2627));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13130 (.out1(R13131), .clock(clock), .in1(_2607));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13131 (.out1(R13132), .clock(clock), .in1(_2596));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13132 (.out1(R13133), .clock(clock), .in1(_2589));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13133 (.out1(R13134), .clock(clock), .in1(_3320));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13134 (.out1(R13135), .clock(clock), .in1(_3225));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13135 (.out1(R13136), .clock(clock), .in1(_3130));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13136 (.out1(R13137), .clock(clock), .in1(_3035));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13137 (.out1(R13138), .clock(clock), .in1(_2940));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13138 (.out1(R13139), .clock(clock), .in1(_2845));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13139 (.out1(R13140), .clock(clock), .in1(_2750));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13140 (.out1(R13141), .clock(clock), .in1(_2655));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13141 (.out1(R13142), .clock(clock), .in1(_2564));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13142 (.out1(R13143), .clock(clock), .in1(_2544));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13143 (.out1(R13144), .clock(clock), .in1(_2535));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13144 (.out1(R13145), .clock(clock), .in1(_2524));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13145 (.out1(R13146), .clock(clock), .in1(_2515));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13146 (.out1(R13147), .clock(clock), .in1(_2504));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13147 (.out1(R13148), .clock(clock), .in1(_2469));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13148 (.out1(R13149), .clock(clock), .in1(_2449));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13149 (.out1(R13150), .clock(clock), .in1(_2440));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13150 (.out1(R13151), .clock(clock), .in1(_2429));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13151 (.out1(R13152), .clock(clock), .in1(_2420));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13152 (.out1(R13153), .clock(clock), .in1(_2409));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13153 (.out1(R13154), .clock(clock), .in1(_2374));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13154 (.out1(R13155), .clock(clock), .in1(_2354));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13155 (.out1(R13156), .clock(clock), .in1(_2345));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13156 (.out1(R13157), .clock(clock), .in1(_2334));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13157 (.out1(R13158), .clock(clock), .in1(_2325));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13158 (.out1(R13159), .clock(clock), .in1(_2314));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13159 (.out1(R13160), .clock(clock), .in1(_2279));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13160 (.out1(R13161), .clock(clock), .in1(_2259));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13161 (.out1(R13162), .clock(clock), .in1(_2250));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13162 (.out1(R13163), .clock(clock), .in1(_2239));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13163 (.out1(R13164), .clock(clock), .in1(_2230));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13164 (.out1(R13165), .clock(clock), .in1(_2219));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13165 (.out1(R13166), .clock(clock), .in1(_2184));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13166 (.out1(R13167), .clock(clock), .in1(_2164));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13167 (.out1(R13168), .clock(clock), .in1(_2155));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13168 (.out1(R13169), .clock(clock), .in1(_2144));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13169 (.out1(R13170), .clock(clock), .in1(_2135));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13170 (.out1(R13171), .clock(clock), .in1(_2124));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13171 (.out1(R13172), .clock(clock), .in1(_2089));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13172 (.out1(R13173), .clock(clock), .in1(_2069));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13173 (.out1(R13174), .clock(clock), .in1(_2060));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13174 (.out1(R13175), .clock(clock), .in1(_2049));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13175 (.out1(R13176), .clock(clock), .in1(_2040));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13176 (.out1(R13177), .clock(clock), .in1(_2029));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13177 (.out1(R13178), .clock(clock), .in1(_1994));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13178 (.out1(R13179), .clock(clock), .in1(_1974));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13179 (.out1(R13180), .clock(clock), .in1(_1965));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13180 (.out1(R13181), .clock(clock), .in1(_1954));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13181 (.out1(R13182), .clock(clock), .in1(_1945));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13182 (.out1(R13183), .clock(clock), .in1(_1934));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13183 (.out1(R13184), .clock(clock), .in1(_1899));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13184 (.out1(R13185), .clock(clock), .in1(_1879));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13185 (.out1(R13186), .clock(clock), .in1(_1870));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13186 (.out1(R13187), .clock(clock), .in1(_1859));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13187 (.out1(R13188), .clock(clock), .in1(_1850));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13188 (.out1(R13189), .clock(clock), .in1(_1839));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13189 (.out1(R13190), .clock(clock), .in1(_1804));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13190 (.out1(R13191), .clock(clock), .in1(_1784));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13191 (.out1(R13192), .clock(clock), .in1(_1775));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13192 (.out1(R13193), .clock(clock), .in1(_1764));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13193 (.out1(R13194), .clock(clock), .in1(_1755));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13194 (.out1(R13195), .clock(clock), .in1(_1744));
  SRAM op3620 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3508),.ADR(R13094));
  SRAM op3613 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3501),.ADR(R13095));
  SRAM op3602 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3490),.ADR(R13096));
  SRAM op3582 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3470),.ADR(R13097));
  SRAM op3522 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3413),.ADR(R13098));
  SRAM op3515 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3406),.ADR(R13099));
  SRAM op3504 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3395),.ADR(R13100));
  SRAM op3484 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3375),.ADR(R13101));
  SRAM op3399 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3293),.ADR(R13102));
  SRAM op3379 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3273),.ADR(R13103));
  SRAM op3368 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3262),.ADR(R13104));
  SRAM op3361 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3255),.ADR(R13105));
  SRAM op3301 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3198),.ADR(R13106));
  SRAM op3281 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3178),.ADR(R13107));
  SRAM op3270 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3167),.ADR(R13108));
  SRAM op3263 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3160),.ADR(R13109));
  SRAM op3203 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3103),.ADR(R13110));
  SRAM op3183 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3083),.ADR(R13111));
  SRAM op3172 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3072),.ADR(R13112));
  SRAM op3165 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3065),.ADR(R13113));
  SRAM op3105 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3008),.ADR(R13114));
  SRAM op3085 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2988),.ADR(R13115));
  SRAM op3074 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2977),.ADR(R13116));
  SRAM op3067 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2970),.ADR(R13117));
  SRAM op3007 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2913),.ADR(R13118));
  SRAM op2987 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2893),.ADR(R13119));
  SRAM op2976 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2882),.ADR(R13120));
  SRAM op2969 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2875),.ADR(R13121));
  SRAM op2909 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2818),.ADR(R13122));
  SRAM op2889 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2798),.ADR(R13123));
  SRAM op2878 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2787),.ADR(R13124));
  SRAM op2871 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2780),.ADR(R13125));
  SRAM op2811 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2723),.ADR(R13126));
  SRAM op2791 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2703),.ADR(R13127));
  SRAM op2780 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2692),.ADR(R13128));
  SRAM op2773 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2685),.ADR(R13129));
  SRAM op2713 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2628),.ADR(R13130));
  SRAM op2693 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2608),.ADR(R13131));
  SRAM op2682 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2597),.ADR(R13132));
  SRAM op2675 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2590),.ADR(R13133));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3427 (.out1(_3321), .in1(R12959), .in2(R13134));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3329 (.out1(_3226), .in1(R12963), .in2(R13135));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3231 (.out1(_3131), .in1(R12967), .in2(R13136));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3133 (.out1(_3036), .in1(R12971), .in2(R13137));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3035 (.out1(_2941), .in1(R12975), .in2(R13138));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2937 (.out1(_2846), .in1(R12979), .in2(R13139));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2839 (.out1(_2751), .in1(R12983), .in2(R13140));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2741 (.out1(_2656), .in1(R12987), .in2(R13141));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2627 (.out1(_2545), .in1(R13143), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2618 (.out1(_2536), .in1(R12991), .in2(R13144));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2587 (.out1(_2505), .in1(R12993), .in2(R13147));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2529 (.out1(_2450), .in1(R13149), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2520 (.out1(_2441), .in1(R12995), .in2(R13150));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2489 (.out1(_2410), .in1(R12997), .in2(R13153));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2431 (.out1(_2355), .in1(R13155), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2422 (.out1(_2346), .in1(R12999), .in2(R13156));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2391 (.out1(_2315), .in1(R13001), .in2(R13159));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2333 (.out1(_2260), .in1(R13161), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2324 (.out1(_2251), .in1(R13003), .in2(R13162));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2293 (.out1(_2220), .in1(R13005), .in2(R13165));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2235 (.out1(_2165), .in1(R13167), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2226 (.out1(_2156), .in1(R13007), .in2(R13168));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2195 (.out1(_2125), .in1(R13009), .in2(R13171));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2137 (.out1(_2070), .in1(R13173), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2128 (.out1(_2061), .in1(R13011), .in2(R13174));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2097 (.out1(_2030), .in1(R13013), .in2(R13177));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2039 (.out1(_1975), .in1(R13179), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2030 (.out1(_1966), .in1(R13015), .in2(R13180));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1999 (.out1(_1935), .in1(R13017), .in2(R13183));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1941 (.out1(_1880), .in1(R13185), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1932 (.out1(_1871), .in1(R13019), .in2(R13186));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1901 (.out1(_1840), .in1(R13021), .in2(R13189));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1843 (.out1(_1785), .in1(R13191), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1834 (.out1(_1776), .in1(R13023), .in2(R13192));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1803 (.out1(_1745), .in1(R13025), .in2(R13195));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op3428 (.out1(_3322), .in1(_3321), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3419 (.out1(_3313), .in1(R13037), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3408 (.out1(_3302), .in1(R13038), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3388 (.out1(_3282), .in1(R13040), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op3330 (.out1(_3227), .in1(_3226), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3321 (.out1(_3218), .in1(R13043), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3310 (.out1(_3207), .in1(R13044), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3290 (.out1(_3187), .in1(R13046), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op3232 (.out1(_3132), .in1(_3131), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3223 (.out1(_3123), .in1(R13049), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3212 (.out1(_3112), .in1(R13050), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3192 (.out1(_3092), .in1(R13052), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op3134 (.out1(_3037), .in1(_3036), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3125 (.out1(_3028), .in1(R13055), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3114 (.out1(_3017), .in1(R13056), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3094 (.out1(_2997), .in1(R13058), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op3036 (.out1(_2942), .in1(_2941), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3027 (.out1(_2933), .in1(R13061), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3016 (.out1(_2922), .in1(R13062), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2996 (.out1(_2902), .in1(R13064), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2938 (.out1(_2847), .in1(_2846), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2929 (.out1(_2838), .in1(R13067), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2918 (.out1(_2827), .in1(R13068), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2898 (.out1(_2807), .in1(R13070), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2840 (.out1(_2752), .in1(_2751), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2831 (.out1(_2743), .in1(R13073), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2820 (.out1(_2732), .in1(R13074), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2800 (.out1(_2712), .in1(R13076), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2742 (.out1(_2657), .in1(_2656), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2733 (.out1(_2648), .in1(R13079), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2722 (.out1(_2637), .in1(R13080), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2702 (.out1(_2617), .in1(R13082), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2647 (.out1(_2565), .in1(R13142), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2628 (.out1(_2546), .in1(_2536), .in2(_2545));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2607 (.out1(_2525), .in1(R13145), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2598 (.out1(_2516), .in1(R12992), .in2(R13146));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2588 (.out1(_2506), .in1(_2505), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2579 (.out1(_2497), .in1(R13085), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2549 (.out1(_2470), .in1(R13148), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2530 (.out1(_2451), .in1(_2441), .in2(_2450));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2509 (.out1(_2430), .in1(R13151), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2500 (.out1(_2421), .in1(R12996), .in2(R13152));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2490 (.out1(_2411), .in1(_2410), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2481 (.out1(_2402), .in1(R13086), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2451 (.out1(_2375), .in1(R13154), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2432 (.out1(_2356), .in1(_2346), .in2(_2355));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2411 (.out1(_2335), .in1(R13157), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2402 (.out1(_2326), .in1(R13000), .in2(R13158));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2392 (.out1(_2316), .in1(_2315), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2383 (.out1(_2307), .in1(R13087), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2353 (.out1(_2280), .in1(R13160), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2334 (.out1(_2261), .in1(_2251), .in2(_2260));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2313 (.out1(_2240), .in1(R13163), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2304 (.out1(_2231), .in1(R13004), .in2(R13164));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2294 (.out1(_2221), .in1(_2220), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2285 (.out1(_2212), .in1(R13088), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2255 (.out1(_2185), .in1(R13166), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2236 (.out1(_2166), .in1(_2156), .in2(_2165));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2215 (.out1(_2145), .in1(R13169), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2206 (.out1(_2136), .in1(R13008), .in2(R13170));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2196 (.out1(_2126), .in1(_2125), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2187 (.out1(_2117), .in1(R13089), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2157 (.out1(_2090), .in1(R13172), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2138 (.out1(_2071), .in1(_2061), .in2(_2070));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2117 (.out1(_2050), .in1(R13175), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2108 (.out1(_2041), .in1(R13012), .in2(R13176));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2098 (.out1(_2031), .in1(_2030), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2089 (.out1(_2022), .in1(R13090), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2059 (.out1(_1995), .in1(R13178), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2040 (.out1(_1976), .in1(_1966), .in2(_1975));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2019 (.out1(_1955), .in1(R13181), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2010 (.out1(_1946), .in1(R13016), .in2(R13182));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2000 (.out1(_1936), .in1(_1935), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1991 (.out1(_1927), .in1(R13091), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1961 (.out1(_1900), .in1(R13184), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1942 (.out1(_1881), .in1(_1871), .in2(_1880));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1921 (.out1(_1860), .in1(R13187), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1912 (.out1(_1851), .in1(R13020), .in2(R13188));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1902 (.out1(_1841), .in1(_1840), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1893 (.out1(_1832), .in1(R13092), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1863 (.out1(_1805), .in1(R13190), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1844 (.out1(_1786), .in1(_1776), .in2(_1785));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1823 (.out1(_1765), .in1(R13193), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1814 (.out1(_1756), .in1(R13024), .in2(R13194));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op1804 (.out1(_1746), .in1(_1745), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1795 (.out1(_1737), .in1(R13093), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2608 (.out1(_2526), .in1(_2516), .in2(_2525));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2510 (.out1(_2431), .in1(_2421), .in2(_2430));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2412 (.out1(_2336), .in1(_2326), .in2(_2335));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2314 (.out1(_2241), .in1(_2231), .in2(_2240));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2216 (.out1(_2146), .in1(_2136), .in2(_2145));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2118 (.out1(_2051), .in1(_2041), .in2(_2050));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2020 (.out1(_1956), .in1(_1946), .in2(_1955));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1922 (.out1(_1861), .in1(_1851), .in2(_1860));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1824 (.out1(_1766), .in1(_1756), .in2(_1765));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3614 (.out1(_3502), .in1(2 'd 2), .in2(R4689));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3603 (.out1(_3491), .in1(2 'd 2), .in2(R4689));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3596 (.out1(_3484), .in1(2 'd 2), .in2(R4689));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3583 (.out1(_3471), .in1(2 'd 2), .in2(R4689));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3576 (.out1(_3464), .in1(2 'd 2), .in2(R4689));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3565 (.out1(_3453), .in1(2 'd 2), .in2(R4689));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3516 (.out1(_3407), .in1(2 'd 2), .in2(R5448));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3505 (.out1(_3396), .in1(2 'd 2), .in2(R5448));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3498 (.out1(_3389), .in1(2 'd 2), .in2(R5448));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3485 (.out1(_3376), .in1(2 'd 2), .in2(R5448));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3478 (.out1(_3369), .in1(2 'd 2), .in2(R5448));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3467 (.out1(_3358), .in1(2 'd 2), .in2(R5448));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3362 (.out1(_3256), .in1(2 'd 2), .in2(R6167));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3264 (.out1(_3161), .in1(2 'd 2), .in2(R6846));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3166 (.out1(_3066), .in1(2 'd 2), .in2(R7485));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3068 (.out1(_2971), .in1(2 'd 2), .in2(R8085));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2970 (.out1(_2876), .in1(2 'd 2), .in2(R8646));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2872 (.out1(_2781), .in1(2 'd 2), .in2(R9168));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2774 (.out1(_2686), .in1(2 'd 2), .in2(R9651));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op2676 (.out1(_2591), .in1(2 'd 2), .in2(R10095));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3594 (.out1(_3482), .in1(leafvec16_3539_D), .in2(R13028));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3574 (.out1(_3462), .in1(leafvec16_3539_D), .in2(R13029));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3563 (.out1(_3451), .in1(leafvec16_3539_D), .in2(R13030));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3556 (.out1(_3444), .in1(leafvec16_3539_D), .in2(R13031));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3496 (.out1(_3387), .in1(leafvec22_3548_D), .in2(R13033));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3476 (.out1(_3367), .in1(leafvec22_3548_D), .in2(R13034));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3465 (.out1(_3356), .in1(leafvec22_3548_D), .in2(R13035));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3458 (.out1(_3349), .in1(leafvec22_3548_D), .in2(R13036));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op3429 (.out1(_3323), .in1(_3322), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3420 (.out1(_3314), .in1(R12960), .in2(_3313));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3409 (.out1(_3303), .in1(R12961), .in2(_3302));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3389 (.out1(_3283), .in1(R12962), .in2(_3282));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op3331 (.out1(_3228), .in1(_3227), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3322 (.out1(_3219), .in1(R12964), .in2(_3218));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3311 (.out1(_3208), .in1(R12965), .in2(_3207));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3291 (.out1(_3188), .in1(R12966), .in2(_3187));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op3233 (.out1(_3133), .in1(_3132), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3224 (.out1(_3124), .in1(R12968), .in2(_3123));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3213 (.out1(_3113), .in1(R12969), .in2(_3112));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3193 (.out1(_3093), .in1(R12970), .in2(_3092));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op3135 (.out1(_3038), .in1(_3037), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3126 (.out1(_3029), .in1(R12972), .in2(_3028));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3115 (.out1(_3018), .in1(R12973), .in2(_3017));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3095 (.out1(_2998), .in1(R12974), .in2(_2997));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op3037 (.out1(_2943), .in1(_2942), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3028 (.out1(_2934), .in1(R12976), .in2(_2933));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3017 (.out1(_2923), .in1(R12977), .in2(_2922));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2997 (.out1(_2903), .in1(R12978), .in2(_2902));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2939 (.out1(_2848), .in1(_2847), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2930 (.out1(_2839), .in1(R12980), .in2(_2838));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2919 (.out1(_2828), .in1(R12981), .in2(_2827));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2899 (.out1(_2808), .in1(R12982), .in2(_2807));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2841 (.out1(_2753), .in1(_2752), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2832 (.out1(_2744), .in1(R12984), .in2(_2743));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2821 (.out1(_2733), .in1(R12985), .in2(_2732));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2801 (.out1(_2713), .in1(R12986), .in2(_2712));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2743 (.out1(_2658), .in1(_2657), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2734 (.out1(_2649), .in1(R12988), .in2(_2648));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2723 (.out1(_2638), .in1(R12989), .in2(_2637));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2703 (.out1(_2618), .in1(R12990), .in2(_2617));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2648 (.out1(_2566), .in1(_2565), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2629 (.out1(_2547), .in1(_2546), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2589 (.out1(_2507), .in1(_2506), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2580 (.out1(_2498), .in1(R12994), .in2(_2497));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2550 (.out1(_2471), .in1(_2470), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2531 (.out1(_2452), .in1(_2451), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2491 (.out1(_2412), .in1(_2411), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2482 (.out1(_2403), .in1(R12998), .in2(_2402));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2452 (.out1(_2376), .in1(_2375), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2433 (.out1(_2357), .in1(_2356), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2393 (.out1(_2317), .in1(_2316), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2384 (.out1(_2308), .in1(R13002), .in2(_2307));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2354 (.out1(_2281), .in1(_2280), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2335 (.out1(_2262), .in1(_2261), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2295 (.out1(_2222), .in1(_2221), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2286 (.out1(_2213), .in1(R13006), .in2(_2212));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2256 (.out1(_2186), .in1(_2185), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2237 (.out1(_2167), .in1(_2166), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2197 (.out1(_2127), .in1(_2126), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2188 (.out1(_2118), .in1(R13010), .in2(_2117));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2158 (.out1(_2091), .in1(_2090), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2139 (.out1(_2072), .in1(_2071), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2099 (.out1(_2032), .in1(_2031), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2090 (.out1(_2023), .in1(R13014), .in2(_2022));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2060 (.out1(_1996), .in1(_1995), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2041 (.out1(_1977), .in1(_1976), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2001 (.out1(_1937), .in1(_1936), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1992 (.out1(_1928), .in1(R13018), .in2(_1927));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1962 (.out1(_1901), .in1(_1900), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1943 (.out1(_1882), .in1(_1881), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1903 (.out1(_1842), .in1(_1841), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1894 (.out1(_1833), .in1(R13022), .in2(_1832));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1864 (.out1(_1806), .in1(_1805), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1845 (.out1(_1787), .in1(_1786), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op1805 (.out1(_1747), .in1(_1746), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1796 (.out1(_1738), .in1(R13026), .in2(_1737));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3622 (.out1(_3510), .in1(R13027), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3524 (.out1(_3415), .in1(R13032), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3430 (.out1(_3324), .in1(_3314), .in2(_3323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op3410 (.out1(_3304), .in1(_3303), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3401 (.out1(_3295), .in1(R13039), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op3390 (.out1(_3284), .in1(_3283), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3381 (.out1(_3275), .in1(R13041), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3370 (.out1(_3264), .in1(R13042), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3332 (.out1(_3229), .in1(_3219), .in2(_3228));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op3312 (.out1(_3209), .in1(_3208), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3303 (.out1(_3200), .in1(R13045), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op3292 (.out1(_3189), .in1(_3188), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3283 (.out1(_3180), .in1(R13047), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3272 (.out1(_3169), .in1(R13048), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3234 (.out1(_3134), .in1(_3124), .in2(_3133));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op3214 (.out1(_3114), .in1(_3113), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3205 (.out1(_3105), .in1(R13051), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op3194 (.out1(_3094), .in1(_3093), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3185 (.out1(_3085), .in1(R13053), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3174 (.out1(_3074), .in1(R13054), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3136 (.out1(_3039), .in1(_3029), .in2(_3038));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op3116 (.out1(_3019), .in1(_3018), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3107 (.out1(_3010), .in1(R13057), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op3096 (.out1(_2999), .in1(_2998), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3087 (.out1(_2990), .in1(R13059), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3076 (.out1(_2979), .in1(R13060), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3038 (.out1(_2944), .in1(_2934), .in2(_2943));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op3018 (.out1(_2924), .in1(_2923), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3009 (.out1(_2915), .in1(R13063), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2998 (.out1(_2904), .in1(_2903), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2989 (.out1(_2895), .in1(R13065), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2978 (.out1(_2884), .in1(R13066), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2940 (.out1(_2849), .in1(_2839), .in2(_2848));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2920 (.out1(_2829), .in1(_2828), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2911 (.out1(_2820), .in1(R13069), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2900 (.out1(_2809), .in1(_2808), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2891 (.out1(_2800), .in1(R13071), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2880 (.out1(_2789), .in1(R13072), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2842 (.out1(_2754), .in1(_2744), .in2(_2753));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2822 (.out1(_2734), .in1(_2733), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2813 (.out1(_2725), .in1(R13075), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2802 (.out1(_2714), .in1(_2713), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2793 (.out1(_2705), .in1(R13077), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2782 (.out1(_2694), .in1(R13078), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2744 (.out1(_2659), .in1(_2649), .in2(_2658));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2724 (.out1(_2639), .in1(_2638), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2715 (.out1(_2630), .in1(R13081), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2704 (.out1(_2619), .in1(_2618), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2695 (.out1(_2610), .in1(R13083), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2684 (.out1(_2599), .in1(R13084), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2649 (.out1(_2567), .in1(_2547), .in2(_2566));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2609 (.out1(_2527), .in1(_2526), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2590 (.out1(_2508), .in1(_2498), .in2(_2507));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2551 (.out1(_2472), .in1(_2452), .in2(_2471));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2511 (.out1(_2432), .in1(_2431), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2492 (.out1(_2413), .in1(_2403), .in2(_2412));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2453 (.out1(_2377), .in1(_2357), .in2(_2376));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2413 (.out1(_2337), .in1(_2336), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2394 (.out1(_2318), .in1(_2308), .in2(_2317));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2355 (.out1(_2282), .in1(_2262), .in2(_2281));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2315 (.out1(_2242), .in1(_2241), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2296 (.out1(_2223), .in1(_2213), .in2(_2222));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2257 (.out1(_2187), .in1(_2167), .in2(_2186));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2217 (.out1(_2147), .in1(_2146), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2198 (.out1(_2128), .in1(_2118), .in2(_2127));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2159 (.out1(_2092), .in1(_2072), .in2(_2091));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2119 (.out1(_2052), .in1(_2051), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2100 (.out1(_2033), .in1(_2023), .in2(_2032));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2061 (.out1(_1997), .in1(_1977), .in2(_1996));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2021 (.out1(_1957), .in1(_1956), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2002 (.out1(_1938), .in1(_1928), .in2(_1937));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1963 (.out1(_1902), .in1(_1882), .in2(_1901));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1923 (.out1(_1862), .in1(_1861), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1904 (.out1(_1843), .in1(_1833), .in2(_1842));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1865 (.out1(_1807), .in1(_1787), .in2(_1806));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1825 (.out1(_1767), .in1(_1766), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1806 (.out1(_1748), .in1(_1738), .in2(_1747));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3933 (.out1(R3934), .clock(clock), .in1(R3933));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4189 (.out1(R4190), .clock(clock), .in1(R4189));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4444 (.out1(R4445), .clock(clock), .in1(R4444));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4689 (.out1(R4690), .clock(clock), .in1(R4689));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4929 (.out1(R4930), .clock(clock), .in1(R4929));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5216 (.out1(R5217), .clock(clock), .in1(R5216));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5448 (.out1(R5449), .clock(clock), .in1(R5448));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5675 (.out1(R5676), .clock(clock), .in1(R5675));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5949 (.out1(R5950), .clock(clock), .in1(R5949));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6380 (.out1(R6381), .clock(clock), .in1(R6380));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6641 (.out1(R6642), .clock(clock), .in1(R6641));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7046 (.out1(R7047), .clock(clock), .in1(R7046));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7293 (.out1(R7294), .clock(clock), .in1(R7293));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7672 (.out1(R7673), .clock(clock), .in1(R7672));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7906 (.out1(R7907), .clock(clock), .in1(R7906));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8259 (.out1(R8260), .clock(clock), .in1(R8259));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8480 (.out1(R8481), .clock(clock), .in1(R8480));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8807 (.out1(R8808), .clock(clock), .in1(R8807));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9015 (.out1(R9016), .clock(clock), .in1(R9015));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9316 (.out1(R9317), .clock(clock), .in1(R9316));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9511 (.out1(R9512), .clock(clock), .in1(R9511));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9786 (.out1(R9787), .clock(clock), .in1(R9786));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9968 (.out1(R9969), .clock(clock), .in1(R9968));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10217 (.out1(R10218), .clock(clock), .in1(R10217));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10386 (.out1(R10387), .clock(clock), .in1(R10386));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10607 (.out1(R10608), .clock(clock), .in1(R10607));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op10763 (.out1(R10764), .clock(clock), .in1(R10763));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10958 (.out1(R10959), .clock(clock), .in1(R10958));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11100 (.out1(R11101), .clock(clock), .in1(R11100));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11269 (.out1(R11270), .clock(clock), .in1(R11269));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11398 (.out1(R11399), .clock(clock), .in1(R11398));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11541 (.out1(R11542), .clock(clock), .in1(R11541));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11657 (.out1(R11658), .clock(clock), .in1(R11657));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11774 (.out1(R11775), .clock(clock), .in1(R11774));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op11877 (.out1(R11878), .clock(clock), .in1(R11877));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11968 (.out1(R11969), .clock(clock), .in1(R11968));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12058 (.out1(R12059), .clock(clock), .in1(R12058));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12123 (.out1(R12124), .clock(clock), .in1(R12123));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12200 (.out1(R12201), .clock(clock), .in1(R12200));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12239 (.out1(R12240), .clock(clock), .in1(R12239));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op12303 (.out1(R12304), .clock(clock), .in1(R12303));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12379 (.out1(R12380), .clock(clock), .in1(R12379));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12390 (.out1(R12391), .clock(clock), .in1(R12390));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12401 (.out1(R12402), .clock(clock), .in1(R12401));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12412 (.out1(R12413), .clock(clock), .in1(R12412));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12423 (.out1(R12424), .clock(clock), .in1(R12423));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12434 (.out1(R12435), .clock(clock), .in1(R12434));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12445 (.out1(R12446), .clock(clock), .in1(R12445));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12456 (.out1(R12457), .clock(clock), .in1(R12456));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12467 (.out1(R12468), .clock(clock), .in1(R12467));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12521 (.out1(R12522), .clock(clock), .in1(R12521));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12532 (.out1(R12533), .clock(clock), .in1(R12532));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12543 (.out1(R12544), .clock(clock), .in1(R12543));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12554 (.out1(R12555), .clock(clock), .in1(R12554));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12565 (.out1(R12566), .clock(clock), .in1(R12565));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12576 (.out1(R12577), .clock(clock), .in1(R12576));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12587 (.out1(R12588), .clock(clock), .in1(R12587));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12598 (.out1(R12599), .clock(clock), .in1(R12598));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12759 (.out1(R12760), .clock(clock), .in1(R12759));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12770 (.out1(R12771), .clock(clock), .in1(R12770));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13195 (.out1(R13196), .clock(clock), .in1(_3508));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13196 (.out1(R13197), .clock(clock), .in1(_3501));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13197 (.out1(R13198), .clock(clock), .in1(_3490));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13198 (.out1(R13199), .clock(clock), .in1(_3470));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13199 (.out1(R13200), .clock(clock), .in1(_3413));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13200 (.out1(R13201), .clock(clock), .in1(_3406));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13201 (.out1(R13202), .clock(clock), .in1(_3395));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13202 (.out1(R13203), .clock(clock), .in1(_3375));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13203 (.out1(R13204), .clock(clock), .in1(_3293));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13204 (.out1(R13205), .clock(clock), .in1(_3273));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13205 (.out1(R13206), .clock(clock), .in1(_3262));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13206 (.out1(R13207), .clock(clock), .in1(_3255));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13207 (.out1(R13208), .clock(clock), .in1(_3198));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13208 (.out1(R13209), .clock(clock), .in1(_3178));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13209 (.out1(R13210), .clock(clock), .in1(_3167));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13210 (.out1(R13211), .clock(clock), .in1(_3160));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13211 (.out1(R13212), .clock(clock), .in1(_3103));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13212 (.out1(R13213), .clock(clock), .in1(_3083));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13213 (.out1(R13214), .clock(clock), .in1(_3072));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13214 (.out1(R13215), .clock(clock), .in1(_3065));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13215 (.out1(R13216), .clock(clock), .in1(_3008));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13216 (.out1(R13217), .clock(clock), .in1(_2988));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13217 (.out1(R13218), .clock(clock), .in1(_2977));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13218 (.out1(R13219), .clock(clock), .in1(_2970));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13219 (.out1(R13220), .clock(clock), .in1(_2913));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13220 (.out1(R13221), .clock(clock), .in1(_2893));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13221 (.out1(R13222), .clock(clock), .in1(_2882));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13222 (.out1(R13223), .clock(clock), .in1(_2875));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13223 (.out1(R13224), .clock(clock), .in1(_2818));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13224 (.out1(R13225), .clock(clock), .in1(_2798));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13225 (.out1(R13226), .clock(clock), .in1(_2787));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13226 (.out1(R13227), .clock(clock), .in1(_2780));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13227 (.out1(R13228), .clock(clock), .in1(_2723));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13228 (.out1(R13229), .clock(clock), .in1(_2703));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13229 (.out1(R13230), .clock(clock), .in1(_2692));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13230 (.out1(R13231), .clock(clock), .in1(_2685));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13231 (.out1(R13232), .clock(clock), .in1(_2628));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13232 (.out1(R13233), .clock(clock), .in1(_2608));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13233 (.out1(R13234), .clock(clock), .in1(_2597));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13234 (.out1(R13235), .clock(clock), .in1(_2590));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13235 (.out1(R13236), .clock(clock), .in1(_3502));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13236 (.out1(R13237), .clock(clock), .in1(_3491));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13237 (.out1(R13238), .clock(clock), .in1(_3484));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13238 (.out1(R13239), .clock(clock), .in1(_3471));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13239 (.out1(R13240), .clock(clock), .in1(_3464));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13240 (.out1(R13241), .clock(clock), .in1(_3453));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13241 (.out1(R13242), .clock(clock), .in1(_3407));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13242 (.out1(R13243), .clock(clock), .in1(_3396));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13243 (.out1(R13244), .clock(clock), .in1(_3389));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13244 (.out1(R13245), .clock(clock), .in1(_3376));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13245 (.out1(R13246), .clock(clock), .in1(_3369));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13246 (.out1(R13247), .clock(clock), .in1(_3358));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13247 (.out1(R13248), .clock(clock), .in1(_3256));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13248 (.out1(R13249), .clock(clock), .in1(_3161));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13249 (.out1(R13250), .clock(clock), .in1(_3066));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13250 (.out1(R13251), .clock(clock), .in1(_2971));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13251 (.out1(R13252), .clock(clock), .in1(_2876));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13252 (.out1(R13253), .clock(clock), .in1(_2781));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13253 (.out1(R13254), .clock(clock), .in1(_2686));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13254 (.out1(R13255), .clock(clock), .in1(_2591));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13255 (.out1(R13256), .clock(clock), .in1(_3482));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13256 (.out1(R13257), .clock(clock), .in1(_3462));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13257 (.out1(R13258), .clock(clock), .in1(_3451));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13258 (.out1(R13259), .clock(clock), .in1(_3444));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13259 (.out1(R13260), .clock(clock), .in1(_3387));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13260 (.out1(R13261), .clock(clock), .in1(_3367));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13261 (.out1(R13262), .clock(clock), .in1(_3356));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13262 (.out1(R13263), .clock(clock), .in1(_3349));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13263 (.out1(R13264), .clock(clock), .in1(_3510));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13264 (.out1(R13265), .clock(clock), .in1(_3415));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13265 (.out1(R13266), .clock(clock), .in1(_3324));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13266 (.out1(R13267), .clock(clock), .in1(_3304));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13267 (.out1(R13268), .clock(clock), .in1(_3295));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13268 (.out1(R13269), .clock(clock), .in1(_3284));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13269 (.out1(R13270), .clock(clock), .in1(_3275));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13270 (.out1(R13271), .clock(clock), .in1(_3264));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13271 (.out1(R13272), .clock(clock), .in1(_3229));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13272 (.out1(R13273), .clock(clock), .in1(_3209));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13273 (.out1(R13274), .clock(clock), .in1(_3200));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13274 (.out1(R13275), .clock(clock), .in1(_3189));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13275 (.out1(R13276), .clock(clock), .in1(_3180));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13276 (.out1(R13277), .clock(clock), .in1(_3169));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13277 (.out1(R13278), .clock(clock), .in1(_3134));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13278 (.out1(R13279), .clock(clock), .in1(_3114));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13279 (.out1(R13280), .clock(clock), .in1(_3105));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13280 (.out1(R13281), .clock(clock), .in1(_3094));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13281 (.out1(R13282), .clock(clock), .in1(_3085));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13282 (.out1(R13283), .clock(clock), .in1(_3074));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13283 (.out1(R13284), .clock(clock), .in1(_3039));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13284 (.out1(R13285), .clock(clock), .in1(_3019));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13285 (.out1(R13286), .clock(clock), .in1(_3010));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13286 (.out1(R13287), .clock(clock), .in1(_2999));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13287 (.out1(R13288), .clock(clock), .in1(_2990));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13288 (.out1(R13289), .clock(clock), .in1(_2979));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13289 (.out1(R13290), .clock(clock), .in1(_2944));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13290 (.out1(R13291), .clock(clock), .in1(_2924));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13291 (.out1(R13292), .clock(clock), .in1(_2915));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13292 (.out1(R13293), .clock(clock), .in1(_2904));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13293 (.out1(R13294), .clock(clock), .in1(_2895));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13294 (.out1(R13295), .clock(clock), .in1(_2884));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13295 (.out1(R13296), .clock(clock), .in1(_2849));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13296 (.out1(R13297), .clock(clock), .in1(_2829));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13297 (.out1(R13298), .clock(clock), .in1(_2820));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13298 (.out1(R13299), .clock(clock), .in1(_2809));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13299 (.out1(R13300), .clock(clock), .in1(_2800));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13300 (.out1(R13301), .clock(clock), .in1(_2789));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13301 (.out1(R13302), .clock(clock), .in1(_2754));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13302 (.out1(R13303), .clock(clock), .in1(_2734));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13303 (.out1(R13304), .clock(clock), .in1(_2725));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13304 (.out1(R13305), .clock(clock), .in1(_2714));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13305 (.out1(R13306), .clock(clock), .in1(_2705));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13306 (.out1(R13307), .clock(clock), .in1(_2694));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13307 (.out1(R13308), .clock(clock), .in1(_2659));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13308 (.out1(R13309), .clock(clock), .in1(_2639));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13309 (.out1(R13310), .clock(clock), .in1(_2630));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13310 (.out1(R13311), .clock(clock), .in1(_2619));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13311 (.out1(R13312), .clock(clock), .in1(_2610));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13312 (.out1(R13313), .clock(clock), .in1(_2599));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13313 (.out1(R13314), .clock(clock), .in1(_2567));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13314 (.out1(R13315), .clock(clock), .in1(_2527));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13315 (.out1(R13316), .clock(clock), .in1(_2508));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13316 (.out1(R13317), .clock(clock), .in1(_2472));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13317 (.out1(R13318), .clock(clock), .in1(_2432));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13318 (.out1(R13319), .clock(clock), .in1(_2413));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13319 (.out1(R13320), .clock(clock), .in1(_2377));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13320 (.out1(R13321), .clock(clock), .in1(_2337));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13321 (.out1(R13322), .clock(clock), .in1(_2318));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13322 (.out1(R13323), .clock(clock), .in1(_2282));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13323 (.out1(R13324), .clock(clock), .in1(_2242));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13324 (.out1(R13325), .clock(clock), .in1(_2223));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13325 (.out1(R13326), .clock(clock), .in1(_2187));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13326 (.out1(R13327), .clock(clock), .in1(_2147));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13327 (.out1(R13328), .clock(clock), .in1(_2128));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13328 (.out1(R13329), .clock(clock), .in1(_2092));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13329 (.out1(R13330), .clock(clock), .in1(_2052));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13330 (.out1(R13331), .clock(clock), .in1(_2033));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13331 (.out1(R13332), .clock(clock), .in1(_1997));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13332 (.out1(R13333), .clock(clock), .in1(_1957));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13333 (.out1(R13334), .clock(clock), .in1(_1938));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13334 (.out1(R13335), .clock(clock), .in1(_1902));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13335 (.out1(R13336), .clock(clock), .in1(_1862));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13336 (.out1(R13337), .clock(clock), .in1(_1843));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13337 (.out1(R13338), .clock(clock), .in1(_1807));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13338 (.out1(R13339), .clock(clock), .in1(_1767));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13339 (.out1(R13340), .clock(clock), .in1(_1748));
  SRAM op3595 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3483),.ADR(R13256));
  SRAM op3575 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3463),.ADR(R13257));
  SRAM op3564 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3452),.ADR(R13258));
  SRAM op3557 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3445),.ADR(R13259));
  SRAM op3497 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3388),.ADR(R13260));
  SRAM op3477 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3368),.ADR(R13261));
  SRAM op3466 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3357),.ADR(R13262));
  SRAM op3459 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3350),.ADR(R13263));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2570 (.out1(_2488), .in1(R10387));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2472 (.out1(_2393), .in1(R10764));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2374 (.out1(_2298), .in1(R11101));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2276 (.out1(_2203), .in1(R11399));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2178 (.out1(_2108), .in1(R11658));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2080 (.out1(_2013), .in1(R11878));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1982 (.out1(_1918), .in1(R12059));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1884 (.out1(_1823), .in1(R12201));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1786 (.out1(_1728), .in1(R12304));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3623 (.out1(_3511), .in1(R13196), .in2(R13264));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3525 (.out1(_3416), .in1(R13200), .in2(R13265));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op3411 (.out1(_3305), .in1(R13267), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3402 (.out1(_3296), .in1(R13204), .in2(R13268));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3371 (.out1(_3265), .in1(R13206), .in2(R13271));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op3313 (.out1(_3210), .in1(R13273), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3304 (.out1(_3201), .in1(R13208), .in2(R13274));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3273 (.out1(_3170), .in1(R13210), .in2(R13277));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op3215 (.out1(_3115), .in1(R13279), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3206 (.out1(_3106), .in1(R13212), .in2(R13280));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3175 (.out1(_3075), .in1(R13214), .in2(R13283));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op3117 (.out1(_3020), .in1(R13285), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3108 (.out1(_3011), .in1(R13216), .in2(R13286));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3077 (.out1(_2980), .in1(R13218), .in2(R13289));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op3019 (.out1(_2925), .in1(R13291), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3010 (.out1(_2916), .in1(R13220), .in2(R13292));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2979 (.out1(_2885), .in1(R13222), .in2(R13295));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2921 (.out1(_2830), .in1(R13297), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2912 (.out1(_2821), .in1(R13224), .in2(R13298));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2881 (.out1(_2790), .in1(R13226), .in2(R13301));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2823 (.out1(_2735), .in1(R13303), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2814 (.out1(_2726), .in1(R13228), .in2(R13304));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2783 (.out1(_2695), .in1(R13230), .in2(R13307));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2725 (.out1(_2640), .in1(R13309), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2716 (.out1(_2631), .in1(R13232), .in2(R13310));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2685 (.out1(_2600), .in1(R13234), .in2(R13313));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2610 (.out1(_2528), .in1(R13315), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2591 (.out1(_2509), .in1(R13316), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2512 (.out1(_2433), .in1(R13318), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2493 (.out1(_2414), .in1(R13319), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2414 (.out1(_2338), .in1(R13321), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2395 (.out1(_2319), .in1(R13322), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2316 (.out1(_2243), .in1(R13324), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2297 (.out1(_2224), .in1(R13325), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2218 (.out1(_2148), .in1(R13327), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2199 (.out1(_2129), .in1(R13328), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2120 (.out1(_2053), .in1(R13330), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2101 (.out1(_2034), .in1(R13331), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2022 (.out1(_1958), .in1(R13333), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2003 (.out1(_1939), .in1(R13334), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1924 (.out1(_1863), .in1(R13336), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1905 (.out1(_1844), .in1(R13337), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1826 (.out1(_1768), .in1(R13339), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op1807 (.out1(_1749), .in1(R13340), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op3624 (.out1(_3512), .in1(_3511), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3615 (.out1(_3503), .in1(R13236), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3604 (.out1(_3492), .in1(R13237), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3584 (.out1(_3472), .in1(R13239), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op3526 (.out1(_3417), .in1(_3416), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3517 (.out1(_3408), .in1(R13242), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3506 (.out1(_3397), .in1(R13243), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3486 (.out1(_3377), .in1(R13245), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3431 (.out1(_3325), .in1(R13266), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3412 (.out1(_3306), .in1(_3296), .in2(_3305));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op3391 (.out1(_3285), .in1(R13269), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3382 (.out1(_3276), .in1(R13205), .in2(R13270));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op3372 (.out1(_3266), .in1(_3265), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3363 (.out1(_3257), .in1(R13248), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3333 (.out1(_3230), .in1(R13272), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3314 (.out1(_3211), .in1(_3201), .in2(_3210));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op3293 (.out1(_3190), .in1(R13275), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3284 (.out1(_3181), .in1(R13209), .in2(R13276));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op3274 (.out1(_3171), .in1(_3170), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3265 (.out1(_3162), .in1(R13249), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3235 (.out1(_3135), .in1(R13278), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3216 (.out1(_3116), .in1(_3106), .in2(_3115));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op3195 (.out1(_3095), .in1(R13281), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3186 (.out1(_3086), .in1(R13213), .in2(R13282));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op3176 (.out1(_3076), .in1(_3075), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3167 (.out1(_3067), .in1(R13250), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3137 (.out1(_3040), .in1(R13284), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3118 (.out1(_3021), .in1(_3011), .in2(_3020));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op3097 (.out1(_3000), .in1(R13287), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3088 (.out1(_2991), .in1(R13217), .in2(R13288));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op3078 (.out1(_2981), .in1(_2980), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3069 (.out1(_2972), .in1(R13251), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3039 (.out1(_2945), .in1(R13290), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3020 (.out1(_2926), .in1(_2916), .in2(_2925));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2999 (.out1(_2905), .in1(R13293), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2990 (.out1(_2896), .in1(R13221), .in2(R13294));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2980 (.out1(_2886), .in1(_2885), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2971 (.out1(_2877), .in1(R13252), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2941 (.out1(_2850), .in1(R13296), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2922 (.out1(_2831), .in1(_2821), .in2(_2830));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2901 (.out1(_2810), .in1(R13299), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2892 (.out1(_2801), .in1(R13225), .in2(R13300));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2882 (.out1(_2791), .in1(_2790), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2873 (.out1(_2782), .in1(R13253), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2843 (.out1(_2755), .in1(R13302), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2824 (.out1(_2736), .in1(_2726), .in2(_2735));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2803 (.out1(_2715), .in1(R13305), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2794 (.out1(_2706), .in1(R13229), .in2(R13306));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2784 (.out1(_2696), .in1(_2695), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2775 (.out1(_2687), .in1(R13254), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2745 (.out1(_2660), .in1(R13308), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2726 (.out1(_2641), .in1(_2631), .in2(_2640));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2705 (.out1(_2620), .in1(R13311), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2696 (.out1(_2611), .in1(R13233), .in2(R13312));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op2686 (.out1(_2601), .in1(_2600), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2677 (.out1(_2592), .in1(R13255), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op2650 (.out1(_2568), .in1(R13314), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2611 (.out1(_2529), .in1(_2509), .in2(_2528));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op2552 (.out1(_2473), .in1(R13317), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2513 (.out1(_2434), .in1(_2414), .in2(_2433));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op2454 (.out1(_2378), .in1(R13320), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2415 (.out1(_2339), .in1(_2319), .in2(_2338));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op2356 (.out1(_2283), .in1(R13323), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2317 (.out1(_2244), .in1(_2224), .in2(_2243));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op2258 (.out1(_2188), .in1(R13326), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2219 (.out1(_2149), .in1(_2129), .in2(_2148));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op2160 (.out1(_2093), .in1(R13329), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2121 (.out1(_2054), .in1(_2034), .in2(_2053));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op2062 (.out1(_1998), .in1(R13332), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2023 (.out1(_1959), .in1(_1939), .in2(_1958));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op1964 (.out1(_1903), .in1(R13335), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1925 (.out1(_1864), .in1(_1844), .in2(_1863));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op1866 (.out1(_1808), .in1(R13338), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1827 (.out1(_1769), .in1(_1749), .in2(_1768));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3392 (.out1(_3286), .in1(_3276), .in2(_3285));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3294 (.out1(_3191), .in1(_3181), .in2(_3190));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3196 (.out1(_3096), .in1(_3086), .in2(_3095));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3098 (.out1(_3001), .in1(_2991), .in2(_3000));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3000 (.out1(_2906), .in1(_2896), .in2(_2905));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2902 (.out1(_2811), .in1(_2801), .in2(_2810));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2804 (.out1(_2716), .in1(_2706), .in2(_2715));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2706 (.out1(_2621), .in1(_2611), .in2(_2620));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3558 (.out1(_3446), .in1(2 'd 2), .in2(R4690));
  LSHIFT_GATE #(.BITSIZE_in1(2), .BITSIZE_in2(32), .BITSIZE_out1(64), .PRECISION(64)) op3460 (.out1(_3351), .in1(2 'd 2), .in2(R5449));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2571 (.out1(_2489), .in1(_2488), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2473 (.out1(_2394), .in1(_2393), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2375 (.out1(_2299), .in1(_2298), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2277 (.out1(_2204), .in1(_2203), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2179 (.out1(_2109), .in1(_2108), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2081 (.out1(_2014), .in1(_2013), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1983 (.out1(_1919), .in1(_1918), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1885 (.out1(_1824), .in1(_1823), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op1787 (.out1(_1729), .in1(_1728), .in2(2 'd 2));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op3625 (.out1(_3513), .in1(_3512), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3616 (.out1(_3504), .in1(R13197), .in2(_3503));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3605 (.out1(_3493), .in1(R13198), .in2(_3492));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3585 (.out1(_3473), .in1(R13199), .in2(_3472));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op3527 (.out1(_3418), .in1(_3417), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3518 (.out1(_3409), .in1(R13201), .in2(_3408));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3507 (.out1(_3398), .in1(R13202), .in2(_3397));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3487 (.out1(_3378), .in1(R13203), .in2(_3377));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op3432 (.out1(_3326), .in1(_3325), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op3413 (.out1(_3307), .in1(_3306), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op3373 (.out1(_3267), .in1(_3266), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3364 (.out1(_3258), .in1(R13207), .in2(_3257));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op3334 (.out1(_3231), .in1(_3230), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op3315 (.out1(_3212), .in1(_3211), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op3275 (.out1(_3172), .in1(_3171), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3266 (.out1(_3163), .in1(R13211), .in2(_3162));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op3236 (.out1(_3136), .in1(_3135), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op3217 (.out1(_3117), .in1(_3116), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op3177 (.out1(_3077), .in1(_3076), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3168 (.out1(_3068), .in1(R13215), .in2(_3067));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op3138 (.out1(_3041), .in1(_3040), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op3119 (.out1(_3022), .in1(_3021), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op3079 (.out1(_2982), .in1(_2981), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3070 (.out1(_2973), .in1(R13219), .in2(_2972));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op3040 (.out1(_2946), .in1(_2945), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op3021 (.out1(_2927), .in1(_2926), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2981 (.out1(_2887), .in1(_2886), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2972 (.out1(_2878), .in1(R13223), .in2(_2877));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2942 (.out1(_2851), .in1(_2850), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2923 (.out1(_2832), .in1(_2831), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2883 (.out1(_2792), .in1(_2791), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2874 (.out1(_2783), .in1(R13227), .in2(_2782));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2844 (.out1(_2756), .in1(_2755), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2825 (.out1(_2737), .in1(_2736), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2785 (.out1(_2697), .in1(_2696), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2776 (.out1(_2688), .in1(R13231), .in2(_2687));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2746 (.out1(_2661), .in1(_2660), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2727 (.out1(_2642), .in1(_2641), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op2687 (.out1(_2602), .in1(_2601), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2678 (.out1(_2593), .in1(R13235), .in2(_2592));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2651 (.out1(_2569), .in1(_2529), .in2(_2568));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2553 (.out1(_2474), .in1(_2434), .in2(_2473));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2455 (.out1(_2379), .in1(_2339), .in2(_2378));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2357 (.out1(_2284), .in1(_2244), .in2(_2283));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2259 (.out1(_2189), .in1(_2149), .in2(_2188));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2161 (.out1(_2094), .in1(_2054), .in2(_2093));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2063 (.out1(_1999), .in1(_1959), .in2(_1998));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1965 (.out1(_1904), .in1(_1864), .in2(_1903));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1867 (.out1(_1809), .in1(_1769), .in2(_1808));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3626 (.out1(_3514), .in1(_3504), .in2(_3513));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op3606 (.out1(_3494), .in1(_3493), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3597 (.out1(_3485), .in1(R13238), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op3586 (.out1(_3474), .in1(_3473), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3577 (.out1(_3465), .in1(R13240), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3566 (.out1(_3454), .in1(R13241), .in2(64 'd 18446744073709551615));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3528 (.out1(_3419), .in1(_3409), .in2(_3418));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op3508 (.out1(_3399), .in1(_3398), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3499 (.out1(_3390), .in1(R13244), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op3488 (.out1(_3379), .in1(_3378), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3479 (.out1(_3370), .in1(R13246), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3468 (.out1(_3359), .in1(R13247), .in2(64 'd 18446744073709551615));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3433 (.out1(_3327), .in1(_3307), .in2(_3326));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3393 (.out1(_3287), .in1(_3286), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3374 (.out1(_3268), .in1(_3258), .in2(_3267));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3335 (.out1(_3232), .in1(_3212), .in2(_3231));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3295 (.out1(_3192), .in1(_3191), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3276 (.out1(_3173), .in1(_3163), .in2(_3172));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3237 (.out1(_3137), .in1(_3117), .in2(_3136));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3197 (.out1(_3097), .in1(_3096), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3178 (.out1(_3078), .in1(_3068), .in2(_3077));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3139 (.out1(_3042), .in1(_3022), .in2(_3041));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3099 (.out1(_3002), .in1(_3001), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3080 (.out1(_2983), .in1(_2973), .in2(_2982));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3041 (.out1(_2947), .in1(_2927), .in2(_2946));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3001 (.out1(_2907), .in1(_2906), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2982 (.out1(_2888), .in1(_2878), .in2(_2887));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2943 (.out1(_2852), .in1(_2832), .in2(_2851));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2903 (.out1(_2812), .in1(_2811), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2884 (.out1(_2793), .in1(_2783), .in2(_2792));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2845 (.out1(_2757), .in1(_2737), .in2(_2756));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2805 (.out1(_2717), .in1(_2716), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2786 (.out1(_2698), .in1(_2688), .in2(_2697));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2747 (.out1(_2662), .in1(_2642), .in2(_2661));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2707 (.out1(_2622), .in1(_2621), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2688 (.out1(_2603), .in1(_2593), .in2(_2602));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op2652 (.out1(_2570), .in1(_2569), .in2(60 'd 1085102592571150095));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op2554 (.out1(_2475), .in1(_2474), .in2(60 'd 1085102592571150095));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op2456 (.out1(_2380), .in1(_2379), .in2(60 'd 1085102592571150095));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op2358 (.out1(_2285), .in1(_2284), .in2(60 'd 1085102592571150095));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op2260 (.out1(_2190), .in1(_2189), .in2(60 'd 1085102592571150095));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op2162 (.out1(_2095), .in1(_2094), .in2(60 'd 1085102592571150095));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op2064 (.out1(_2000), .in1(_1999), .in2(60 'd 1085102592571150095));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op1966 (.out1(_1905), .in1(_1904), .in2(60 'd 1085102592571150095));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op1868 (.out1(_1810), .in1(_1809), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3934 (.out1(R3935), .clock(clock), .in1(R3934));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4190 (.out1(R4191), .clock(clock), .in1(R4190));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4445 (.out1(R4446), .clock(clock), .in1(R4445));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4930 (.out1(R4931), .clock(clock), .in1(R4930));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5217 (.out1(R5218), .clock(clock), .in1(R5217));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5676 (.out1(R5677), .clock(clock), .in1(R5676));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5950 (.out1(R5951), .clock(clock), .in1(R5950));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6381 (.out1(R6382), .clock(clock), .in1(R6381));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op6642 (.out1(R6643), .clock(clock), .in1(R6642));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7047 (.out1(R7048), .clock(clock), .in1(R7047));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7294 (.out1(R7295), .clock(clock), .in1(R7294));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7673 (.out1(R7674), .clock(clock), .in1(R7673));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op7907 (.out1(R7908), .clock(clock), .in1(R7907));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8260 (.out1(R8261), .clock(clock), .in1(R8260));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op8481 (.out1(R8482), .clock(clock), .in1(R8481));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8808 (.out1(R8809), .clock(clock), .in1(R8808));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9016 (.out1(R9017), .clock(clock), .in1(R9016));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9317 (.out1(R9318), .clock(clock), .in1(R9317));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9512 (.out1(R9513), .clock(clock), .in1(R9512));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9787 (.out1(R9788), .clock(clock), .in1(R9787));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op9969 (.out1(R9970), .clock(clock), .in1(R9969));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10218 (.out1(R10219), .clock(clock), .in1(R10218));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10608 (.out1(R10609), .clock(clock), .in1(R10608));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10959 (.out1(R10960), .clock(clock), .in1(R10959));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11270 (.out1(R11271), .clock(clock), .in1(R11270));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11542 (.out1(R11543), .clock(clock), .in1(R11542));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11775 (.out1(R11776), .clock(clock), .in1(R11775));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11969 (.out1(R11970), .clock(clock), .in1(R11969));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12124 (.out1(R12125), .clock(clock), .in1(R12124));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12240 (.out1(R12241), .clock(clock), .in1(R12240));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12380 (.out1(R12381), .clock(clock), .in1(R12380));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12391 (.out1(R12392), .clock(clock), .in1(R12391));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12402 (.out1(R12403), .clock(clock), .in1(R12402));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12413 (.out1(R12414), .clock(clock), .in1(R12413));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12424 (.out1(R12425), .clock(clock), .in1(R12424));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12435 (.out1(R12436), .clock(clock), .in1(R12435));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12446 (.out1(R12447), .clock(clock), .in1(R12446));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12457 (.out1(R12458), .clock(clock), .in1(R12457));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12468 (.out1(R12469), .clock(clock), .in1(R12468));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12522 (.out1(R12523), .clock(clock), .in1(R12522));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12533 (.out1(R12534), .clock(clock), .in1(R12533));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12544 (.out1(R12545), .clock(clock), .in1(R12544));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12555 (.out1(R12556), .clock(clock), .in1(R12555));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12566 (.out1(R12567), .clock(clock), .in1(R12566));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12577 (.out1(R12578), .clock(clock), .in1(R12577));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12588 (.out1(R12589), .clock(clock), .in1(R12588));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12599 (.out1(R12600), .clock(clock), .in1(R12599));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12760 (.out1(R12761), .clock(clock), .in1(R12760));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12771 (.out1(R12772), .clock(clock), .in1(R12771));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13340 (.out1(R13341), .clock(clock), .in1(_3483));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13341 (.out1(R13342), .clock(clock), .in1(_3463));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13342 (.out1(R13343), .clock(clock), .in1(_3452));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13343 (.out1(R13344), .clock(clock), .in1(_3445));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13344 (.out1(R13345), .clock(clock), .in1(_3388));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13345 (.out1(R13346), .clock(clock), .in1(_3368));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13346 (.out1(R13347), .clock(clock), .in1(_3357));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13347 (.out1(R13348), .clock(clock), .in1(_3350));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13348 (.out1(R13349), .clock(clock), .in1(_3446));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13349 (.out1(R13350), .clock(clock), .in1(_3351));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13350 (.out1(R13351), .clock(clock), .in1(_2489));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13351 (.out1(R13352), .clock(clock), .in1(_2394));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13352 (.out1(R13353), .clock(clock), .in1(_2299));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13353 (.out1(R13354), .clock(clock), .in1(_2204));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13354 (.out1(R13355), .clock(clock), .in1(_2109));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13355 (.out1(R13356), .clock(clock), .in1(_2014));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13356 (.out1(R13357), .clock(clock), .in1(_1919));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13357 (.out1(R13358), .clock(clock), .in1(_1824));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13358 (.out1(R13359), .clock(clock), .in1(_1729));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13359 (.out1(R13360), .clock(clock), .in1(_3514));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13360 (.out1(R13361), .clock(clock), .in1(_3494));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13361 (.out1(R13362), .clock(clock), .in1(_3485));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13362 (.out1(R13363), .clock(clock), .in1(_3474));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13363 (.out1(R13364), .clock(clock), .in1(_3465));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13364 (.out1(R13365), .clock(clock), .in1(_3454));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13365 (.out1(R13366), .clock(clock), .in1(_3419));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13366 (.out1(R13367), .clock(clock), .in1(_3399));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13367 (.out1(R13368), .clock(clock), .in1(_3390));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13368 (.out1(R13369), .clock(clock), .in1(_3379));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13369 (.out1(R13370), .clock(clock), .in1(_3370));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13370 (.out1(R13371), .clock(clock), .in1(_3359));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13371 (.out1(R13372), .clock(clock), .in1(_3327));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13372 (.out1(R13373), .clock(clock), .in1(_3287));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13373 (.out1(R13374), .clock(clock), .in1(_3268));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13374 (.out1(R13375), .clock(clock), .in1(_3232));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13375 (.out1(R13376), .clock(clock), .in1(_3192));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13376 (.out1(R13377), .clock(clock), .in1(_3173));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13377 (.out1(R13378), .clock(clock), .in1(_3137));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13378 (.out1(R13379), .clock(clock), .in1(_3097));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13379 (.out1(R13380), .clock(clock), .in1(_3078));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13380 (.out1(R13381), .clock(clock), .in1(_3042));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13381 (.out1(R13382), .clock(clock), .in1(_3002));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13382 (.out1(R13383), .clock(clock), .in1(_2983));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13383 (.out1(R13384), .clock(clock), .in1(_2947));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13384 (.out1(R13385), .clock(clock), .in1(_2907));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13385 (.out1(R13386), .clock(clock), .in1(_2888));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13386 (.out1(R13387), .clock(clock), .in1(_2852));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13387 (.out1(R13388), .clock(clock), .in1(_2812));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13388 (.out1(R13389), .clock(clock), .in1(_2793));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13389 (.out1(R13390), .clock(clock), .in1(_2757));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13390 (.out1(R13391), .clock(clock), .in1(_2717));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13391 (.out1(R13392), .clock(clock), .in1(_2698));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13392 (.out1(R13393), .clock(clock), .in1(_2662));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13393 (.out1(R13394), .clock(clock), .in1(_2622));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13394 (.out1(R13395), .clock(clock), .in1(_2603));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13395 (.out1(R13396), .clock(clock), .in1(_2570));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13396 (.out1(R13397), .clock(clock), .in1(_2475));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13397 (.out1(R13398), .clock(clock), .in1(_2380));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13398 (.out1(R13399), .clock(clock), .in1(_2285));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13399 (.out1(R13400), .clock(clock), .in1(_2190));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13400 (.out1(R13401), .clock(clock), .in1(_2095));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13401 (.out1(R13402), .clock(clock), .in1(_2000));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13402 (.out1(R13403), .clock(clock), .in1(_1905));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13403 (.out1(R13404), .clock(clock), .in1(_1810));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op2653 (.out1(_2571), .in1(R13396), .in2(57 'd 72340172838076673));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op2555 (.out1(_2476), .in1(R13397), .in2(57 'd 72340172838076673));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op2457 (.out1(_2381), .in1(R13398), .in2(57 'd 72340172838076673));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op2359 (.out1(_2286), .in1(R13399), .in2(57 'd 72340172838076673));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op2261 (.out1(_2191), .in1(R13400), .in2(57 'd 72340172838076673));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op2163 (.out1(_2096), .in1(R13401), .in2(57 'd 72340172838076673));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op2065 (.out1(_2001), .in1(R13402), .in2(57 'd 72340172838076673));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op1967 (.out1(_1906), .in1(R13403), .in2(57 'd 72340172838076673));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op1869 (.out1(_1811), .in1(R13404), .in2(57 'd 72340172838076673));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3354 (.out1(_3248), .in1(R5951));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3256 (.out1(_3153), .in1(R6643));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3158 (.out1(_3058), .in1(R7295));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3060 (.out1(_2963), .in1(R7908));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2962 (.out1(_2868), .in1(R8482));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2864 (.out1(_2773), .in1(R9017));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2766 (.out1(_2678), .in1(R9513));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2668 (.out1(_2583), .in1(R9970));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op3607 (.out1(_3495), .in1(R13361), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3598 (.out1(_3486), .in1(R13341), .in2(R13362));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3567 (.out1(_3455), .in1(R13343), .in2(R13365));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op3509 (.out1(_3400), .in1(R13367), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3500 (.out1(_3391), .in1(R13345), .in2(R13368));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3469 (.out1(_3360), .in1(R13347), .in2(R13371));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op3394 (.out1(_3288), .in1(R13373), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op3375 (.out1(_3269), .in1(R13374), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op3296 (.out1(_3193), .in1(R13376), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op3277 (.out1(_3174), .in1(R13377), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op3198 (.out1(_3098), .in1(R13379), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op3179 (.out1(_3079), .in1(R13380), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op3100 (.out1(_3003), .in1(R13382), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op3081 (.out1(_2984), .in1(R13383), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op3002 (.out1(_2908), .in1(R13385), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2983 (.out1(_2889), .in1(R13386), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2904 (.out1(_2813), .in1(R13388), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2885 (.out1(_2794), .in1(R13389), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2806 (.out1(_2718), .in1(R13391), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2787 (.out1(_2699), .in1(R13392), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2708 (.out1(_2623), .in1(R13394), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op2689 (.out1(_2604), .in1(R13395), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3627 (.out1(_3515), .in1(R13360), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3608 (.out1(_3496), .in1(_3486), .in2(_3495));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op3587 (.out1(_3475), .in1(R13363), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3578 (.out1(_3466), .in1(R13342), .in2(R13364));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op3568 (.out1(_3456), .in1(_3455), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3559 (.out1(_3447), .in1(R13349), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3529 (.out1(_3420), .in1(R13366), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3510 (.out1(_3401), .in1(_3391), .in2(_3400));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op3489 (.out1(_3380), .in1(R13369), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3480 (.out1(_3371), .in1(R13346), .in2(R13370));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(1), .BITSIZE_out1(64), .PRECISION(64)) op3470 (.out1(_3361), .in1(_3360), .in2(1 'd 1));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3461 (.out1(_3352), .in1(R13350), .in2(64 'd 18446744073709551615));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op3434 (.out1(_3328), .in1(R13372), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3395 (.out1(_3289), .in1(_3269), .in2(_3288));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op3336 (.out1(_3233), .in1(R13375), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3297 (.out1(_3194), .in1(_3174), .in2(_3193));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op3238 (.out1(_3138), .in1(R13378), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3199 (.out1(_3099), .in1(_3079), .in2(_3098));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op3140 (.out1(_3043), .in1(R13381), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3101 (.out1(_3004), .in1(_2984), .in2(_3003));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op3042 (.out1(_2948), .in1(R13384), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3003 (.out1(_2909), .in1(_2889), .in2(_2908));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op2944 (.out1(_2853), .in1(R13387), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2905 (.out1(_2814), .in1(_2794), .in2(_2813));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op2846 (.out1(_2758), .in1(R13390), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2807 (.out1(_2719), .in1(_2699), .in2(_2718));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op2748 (.out1(_2663), .in1(R13393), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2709 (.out1(_2624), .in1(_2604), .in2(_2623));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3588 (.out1(_3476), .in1(_3466), .in2(_3475));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3490 (.out1(_3381), .in1(_3371), .in2(_3380));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3355 (.out1(_3249), .in1(_3248), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3257 (.out1(_3154), .in1(_3153), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3159 (.out1(_3059), .in1(_3058), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3061 (.out1(_2964), .in1(_2963), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2963 (.out1(_2869), .in1(_2868), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2865 (.out1(_2774), .in1(_2773), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2767 (.out1(_2679), .in1(_2678), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op2669 (.out1(_2584), .in1(_2583), .in2(2 'd 2));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2572 (.out1(_2490), .in1(base1_76_3622_D), .in2(R13351));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2474 (.out1(_2395), .in1(base1_82_3630_D), .in2(R13352));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2376 (.out1(_2300), .in1(base1_88_3638_D), .in2(R13353));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2278 (.out1(_2205), .in1(base1_94_3646_D), .in2(R13354));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2180 (.out1(_2110), .in1(base1_100_3654_D), .in2(R13355));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2082 (.out1(_2015), .in1(base1_106_3662_D), .in2(R13356));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1984 (.out1(_1920), .in1(base1_112_3670_D), .in2(R13357));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1886 (.out1(_1825), .in1(base1_118_3678_D), .in2(R13358));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1788 (.out1(_1730), .in1(base1_124_3685_D), .in2(R13359));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op3628 (.out1(_3516), .in1(_3515), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op3609 (.out1(_3497), .in1(_3496), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op3569 (.out1(_3457), .in1(_3456), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3560 (.out1(_3448), .in1(R13344), .in2(_3447));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op3530 (.out1(_3421), .in1(_3420), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op3511 (.out1(_3402), .in1(_3401), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(63), .BITSIZE_out1(64)) op3471 (.out1(_3362), .in1(_3361), .in2(63 'd 6148914691236517205));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3462 (.out1(_3353), .in1(R13348), .in2(_3352));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3435 (.out1(_3329), .in1(_3289), .in2(_3328));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3337 (.out1(_3234), .in1(_3194), .in2(_3233));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3239 (.out1(_3139), .in1(_3099), .in2(_3138));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3141 (.out1(_3044), .in1(_3004), .in2(_3043));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3043 (.out1(_2949), .in1(_2909), .in2(_2948));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2945 (.out1(_2854), .in1(_2814), .in2(_2853));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2847 (.out1(_2759), .in1(_2719), .in2(_2758));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2749 (.out1(_2664), .in1(_2624), .in2(_2663));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3629 (.out1(_3517), .in1(_3497), .in2(_3516));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3589 (.out1(_3477), .in1(_3476), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3570 (.out1(_3458), .in1(_3448), .in2(_3457));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3531 (.out1(_3422), .in1(_3402), .in2(_3421));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3491 (.out1(_3382), .in1(_3381), .in2(2 'd 2));
  SUB_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3472 (.out1(_3363), .in1(_3353), .in2(_3362));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op3436 (.out1(_3330), .in1(_3329), .in2(60 'd 1085102592571150095));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op3338 (.out1(_3235), .in1(_3234), .in2(60 'd 1085102592571150095));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op3240 (.out1(_3140), .in1(_3139), .in2(60 'd 1085102592571150095));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op3142 (.out1(_3045), .in1(_3044), .in2(60 'd 1085102592571150095));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op3044 (.out1(_2950), .in1(_2949), .in2(60 'd 1085102592571150095));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op2946 (.out1(_2855), .in1(_2854), .in2(60 'd 1085102592571150095));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op2848 (.out1(_2760), .in1(_2759), .in2(60 'd 1085102592571150095));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op2750 (.out1(_2665), .in1(_2664), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3935 (.out1(R3936), .clock(clock), .in1(R3935));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4191 (.out1(R4192), .clock(clock), .in1(R4191));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op4446 (.out1(R4447), .clock(clock), .in1(R4446));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4931 (.out1(R4932), .clock(clock), .in1(R4931));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op5218 (.out1(R5219), .clock(clock), .in1(R5218));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5677 (.out1(R5678), .clock(clock), .in1(R5677));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6382 (.out1(R6383), .clock(clock), .in1(R6382));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7048 (.out1(R7049), .clock(clock), .in1(R7048));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7674 (.out1(R7675), .clock(clock), .in1(R7674));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8261 (.out1(R8262), .clock(clock), .in1(R8261));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8809 (.out1(R8810), .clock(clock), .in1(R8809));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9318 (.out1(R9319), .clock(clock), .in1(R9318));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9788 (.out1(R9789), .clock(clock), .in1(R9788));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10219 (.out1(R10220), .clock(clock), .in1(R10219));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10609 (.out1(R10610), .clock(clock), .in1(R10609));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10960 (.out1(R10961), .clock(clock), .in1(R10960));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11271 (.out1(R11272), .clock(clock), .in1(R11271));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11543 (.out1(R11544), .clock(clock), .in1(R11543));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11776 (.out1(R11777), .clock(clock), .in1(R11776));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11970 (.out1(R11971), .clock(clock), .in1(R11970));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12125 (.out1(R12126), .clock(clock), .in1(R12125));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12241 (.out1(R12242), .clock(clock), .in1(R12241));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12381 (.out1(R12382), .clock(clock), .in1(R12381));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12392 (.out1(R12393), .clock(clock), .in1(R12392));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12403 (.out1(R12404), .clock(clock), .in1(R12403));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12414 (.out1(R12415), .clock(clock), .in1(R12414));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12425 (.out1(R12426), .clock(clock), .in1(R12425));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12436 (.out1(R12437), .clock(clock), .in1(R12436));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12447 (.out1(R12448), .clock(clock), .in1(R12447));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12458 (.out1(R12459), .clock(clock), .in1(R12458));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12469 (.out1(R12470), .clock(clock), .in1(R12469));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12523 (.out1(R12524), .clock(clock), .in1(R12523));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12534 (.out1(R12535), .clock(clock), .in1(R12534));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12545 (.out1(R12546), .clock(clock), .in1(R12545));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12556 (.out1(R12557), .clock(clock), .in1(R12556));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12567 (.out1(R12568), .clock(clock), .in1(R12567));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12578 (.out1(R12579), .clock(clock), .in1(R12578));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12589 (.out1(R12590), .clock(clock), .in1(R12589));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12600 (.out1(R12601), .clock(clock), .in1(R12600));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12761 (.out1(R12762), .clock(clock), .in1(R12761));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12772 (.out1(R12773), .clock(clock), .in1(R12772));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13404 (.out1(R13405), .clock(clock), .in1(_2571));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13405 (.out1(R13406), .clock(clock), .in1(_2476));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13406 (.out1(R13407), .clock(clock), .in1(_2381));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13407 (.out1(R13408), .clock(clock), .in1(_2286));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13408 (.out1(R13409), .clock(clock), .in1(_2191));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13409 (.out1(R13410), .clock(clock), .in1(_2096));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13410 (.out1(R13411), .clock(clock), .in1(_2001));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13411 (.out1(R13412), .clock(clock), .in1(_1906));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13412 (.out1(R13413), .clock(clock), .in1(_1811));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13413 (.out1(R13414), .clock(clock), .in1(_3249));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13414 (.out1(R13415), .clock(clock), .in1(_3154));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13415 (.out1(R13416), .clock(clock), .in1(_3059));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13416 (.out1(R13417), .clock(clock), .in1(_2964));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13417 (.out1(R13418), .clock(clock), .in1(_2869));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13418 (.out1(R13419), .clock(clock), .in1(_2774));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13419 (.out1(R13420), .clock(clock), .in1(_2679));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13420 (.out1(R13421), .clock(clock), .in1(_2584));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13421 (.out1(R13422), .clock(clock), .in1(_2490));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13422 (.out1(R13423), .clock(clock), .in1(_2395));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13423 (.out1(R13424), .clock(clock), .in1(_2300));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13424 (.out1(R13425), .clock(clock), .in1(_2205));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13425 (.out1(R13426), .clock(clock), .in1(_2110));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13426 (.out1(R13427), .clock(clock), .in1(_2015));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13427 (.out1(R13428), .clock(clock), .in1(_1920));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13428 (.out1(R13429), .clock(clock), .in1(_1825));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13429 (.out1(R13430), .clock(clock), .in1(_1730));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13430 (.out1(R13431), .clock(clock), .in1(_3517));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13431 (.out1(R13432), .clock(clock), .in1(_3477));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13432 (.out1(R13433), .clock(clock), .in1(_3458));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13433 (.out1(R13434), .clock(clock), .in1(_3422));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13434 (.out1(R13435), .clock(clock), .in1(_3382));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13435 (.out1(R13436), .clock(clock), .in1(_3363));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13436 (.out1(R13437), .clock(clock), .in1(_3330));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13437 (.out1(R13438), .clock(clock), .in1(_3235));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13438 (.out1(R13439), .clock(clock), .in1(_3140));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13439 (.out1(R13440), .clock(clock), .in1(_3045));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13440 (.out1(R13441), .clock(clock), .in1(_2950));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13441 (.out1(R13442), .clock(clock), .in1(_2855));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13442 (.out1(R13443), .clock(clock), .in1(_2760));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13443 (.out1(R13444), .clock(clock), .in1(_2665));
  SRAM op2573 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2491),.ADR(R13422));
  SRAM op2475 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2396),.ADR(R13423));
  SRAM op2377 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2301),.ADR(R13424));
  SRAM op2279 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2206),.ADR(R13425));
  SRAM op2181 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2111),.ADR(R13426));
  SRAM op2083 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2016),.ADR(R13427));
  SRAM op1985 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1921),.ADR(R13428));
  SRAM op1887 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1826),.ADR(R13429));
  SRAM op1789 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_1731),.ADR(R13430));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op3437 (.out1(_3331), .in1(R13437), .in2(57 'd 72340172838076673));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op3339 (.out1(_3236), .in1(R13438), .in2(57 'd 72340172838076673));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op3241 (.out1(_3141), .in1(R13439), .in2(57 'd 72340172838076673));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op3143 (.out1(_3046), .in1(R13440), .in2(57 'd 72340172838076673));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op3045 (.out1(_2951), .in1(R13441), .in2(57 'd 72340172838076673));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op2947 (.out1(_2856), .in1(R13442), .in2(57 'd 72340172838076673));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op2849 (.out1(_2761), .in1(R13443), .in2(57 'd 72340172838076673));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op2751 (.out1(_2666), .in1(R13444), .in2(57 'd 72340172838076673));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3550 (.out1(_3438), .in1(R4447));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3452 (.out1(_3343), .in1(R5219));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op3590 (.out1(_3478), .in1(R13432), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op3571 (.out1(_3459), .in1(R13433), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op3492 (.out1(_3383), .in1(R13435), .in2(62 'd 3689348814741910323));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(62), .BITSIZE_out1(64)) op3473 (.out1(_3364), .in1(R13436), .in2(62 'd 3689348814741910323));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op3630 (.out1(_3518), .in1(R13431), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3591 (.out1(_3479), .in1(_3459), .in2(_3478));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(3), .BITSIZE_out1(64), .PRECISION(64)) op3532 (.out1(_3423), .in1(R13434), .in2(3 'd 4));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3493 (.out1(_3384), .in1(_3364), .in2(_3383));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3551 (.out1(_3439), .in1(_3438), .in2(2 'd 2));
  LSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(2), .BITSIZE_out1(64), .PRECISION(64)) op3453 (.out1(_3344), .in1(_3343), .in2(2 'd 2));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3356 (.out1(_3250), .in1(base1_28_3557_D), .in2(R13414));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3258 (.out1(_3155), .in1(base1_34_3565_D), .in2(R13415));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3160 (.out1(_3060), .in1(base1_40_3573_D), .in2(R13416));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3062 (.out1(_2965), .in1(base1_46_3581_D), .in2(R13417));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2964 (.out1(_2870), .in1(base1_52_3589_D), .in2(R13418));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2866 (.out1(_2775), .in1(base1_58_3597_D), .in2(R13419));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2768 (.out1(_2680), .in1(base1_64_3606_D), .in2(R13420));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2670 (.out1(_2585), .in1(base1_70_3614_D), .in2(R13421));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3631 (.out1(_3519), .in1(_3479), .in2(_3518));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3533 (.out1(_3424), .in1(_3384), .in2(_3423));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op2654 (.out1(_2572), .in1(R13405), .in2(6 'd 56));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op2556 (.out1(_2477), .in1(R13406), .in2(6 'd 56));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op2458 (.out1(_2382), .in1(R13407), .in2(6 'd 56));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op2360 (.out1(_2287), .in1(R13408), .in2(6 'd 56));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op2262 (.out1(_2192), .in1(R13409), .in2(6 'd 56));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op2164 (.out1(_2097), .in1(R13410), .in2(6 'd 56));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op2066 (.out1(_2002), .in1(R13411), .in2(6 'd 56));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op1968 (.out1(_1907), .in1(R13412), .in2(6 'd 56));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op1870 (.out1(_1812), .in1(R13413), .in2(6 'd 56));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op3632 (.out1(_3520), .in1(_3519), .in2(60 'd 1085102592571150095));
  bit_and #(.BITSIZE_in1(64), .BITSIZE_in2(60), .BITSIZE_out1(64)) op3534 (.out1(_3425), .in1(_3424), .in2(60 'd 1085102592571150095));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3936 (.out1(R3937), .clock(clock), .in1(R3936));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4192 (.out1(R4193), .clock(clock), .in1(R4192));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4932 (.out1(R4933), .clock(clock), .in1(R4932));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5678 (.out1(R5679), .clock(clock), .in1(R5678));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6383 (.out1(R6384), .clock(clock), .in1(R6383));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7049 (.out1(R7050), .clock(clock), .in1(R7049));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7675 (.out1(R7676), .clock(clock), .in1(R7675));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8262 (.out1(R8263), .clock(clock), .in1(R8262));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8810 (.out1(R8811), .clock(clock), .in1(R8810));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9319 (.out1(R9320), .clock(clock), .in1(R9319));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9789 (.out1(R9790), .clock(clock), .in1(R9789));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10220 (.out1(R10221), .clock(clock), .in1(R10220));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10610 (.out1(R10611), .clock(clock), .in1(R10610));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10961 (.out1(R10962), .clock(clock), .in1(R10961));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11272 (.out1(R11273), .clock(clock), .in1(R11272));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11544 (.out1(R11545), .clock(clock), .in1(R11544));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11777 (.out1(R11778), .clock(clock), .in1(R11777));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11971 (.out1(R11972), .clock(clock), .in1(R11971));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12126 (.out1(R12127), .clock(clock), .in1(R12126));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12242 (.out1(R12243), .clock(clock), .in1(R12242));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12382 (.out1(R12383), .clock(clock), .in1(R12382));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12393 (.out1(R12394), .clock(clock), .in1(R12393));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12404 (.out1(R12405), .clock(clock), .in1(R12404));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12415 (.out1(R12416), .clock(clock), .in1(R12415));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12426 (.out1(R12427), .clock(clock), .in1(R12426));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12437 (.out1(R12438), .clock(clock), .in1(R12437));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12448 (.out1(R12449), .clock(clock), .in1(R12448));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12459 (.out1(R12460), .clock(clock), .in1(R12459));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12470 (.out1(R12471), .clock(clock), .in1(R12470));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12524 (.out1(R12525), .clock(clock), .in1(R12524));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12535 (.out1(R12536), .clock(clock), .in1(R12535));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12546 (.out1(R12547), .clock(clock), .in1(R12546));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12557 (.out1(R12558), .clock(clock), .in1(R12557));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12568 (.out1(R12569), .clock(clock), .in1(R12568));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12579 (.out1(R12580), .clock(clock), .in1(R12579));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12590 (.out1(R12591), .clock(clock), .in1(R12590));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12601 (.out1(R12602), .clock(clock), .in1(R12601));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12762 (.out1(R12763), .clock(clock), .in1(R12762));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12773 (.out1(R12774), .clock(clock), .in1(R12773));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13444 (.out1(R13445), .clock(clock), .in1(_2491));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13445 (.out1(R13446), .clock(clock), .in1(_2396));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13446 (.out1(R13447), .clock(clock), .in1(_2301));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13447 (.out1(R13448), .clock(clock), .in1(_2206));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13448 (.out1(R13449), .clock(clock), .in1(_2111));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13449 (.out1(R13450), .clock(clock), .in1(_2016));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13450 (.out1(R13451), .clock(clock), .in1(_1921));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13451 (.out1(R13452), .clock(clock), .in1(_1826));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13452 (.out1(R13453), .clock(clock), .in1(_1731));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13453 (.out1(R13454), .clock(clock), .in1(_3331));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13454 (.out1(R13455), .clock(clock), .in1(_3236));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13455 (.out1(R13456), .clock(clock), .in1(_3141));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13456 (.out1(R13457), .clock(clock), .in1(_3046));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13457 (.out1(R13458), .clock(clock), .in1(_2951));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13458 (.out1(R13459), .clock(clock), .in1(_2856));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13459 (.out1(R13460), .clock(clock), .in1(_2761));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13460 (.out1(R13461), .clock(clock), .in1(_2666));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13461 (.out1(R13462), .clock(clock), .in1(_3439));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13462 (.out1(R13463), .clock(clock), .in1(_3344));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13463 (.out1(R13464), .clock(clock), .in1(_3250));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13464 (.out1(R13465), .clock(clock), .in1(_3155));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13465 (.out1(R13466), .clock(clock), .in1(_3060));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13466 (.out1(R13467), .clock(clock), .in1(_2965));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13467 (.out1(R13468), .clock(clock), .in1(_2870));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13468 (.out1(R13469), .clock(clock), .in1(_2775));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13469 (.out1(R13470), .clock(clock), .in1(_2680));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13470 (.out1(R13471), .clock(clock), .in1(_2585));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13471 (.out1(R13472), .clock(clock), .in1(_2572));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13472 (.out1(R13473), .clock(clock), .in1(_2477));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13473 (.out1(R13474), .clock(clock), .in1(_2382));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13474 (.out1(R13475), .clock(clock), .in1(_2287));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13475 (.out1(R13476), .clock(clock), .in1(_2192));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13476 (.out1(R13477), .clock(clock), .in1(_2097));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13477 (.out1(R13478), .clock(clock), .in1(_2002));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13478 (.out1(R13479), .clock(clock), .in1(_1907));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13479 (.out1(R13480), .clock(clock), .in1(_1812));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13480 (.out1(R13481), .clock(clock), .in1(_3520));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13481 (.out1(R13482), .clock(clock), .in1(_3425));
  SRAM op3357 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3251),.ADR(R13464));
  SRAM op3259 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3156),.ADR(R13465));
  SRAM op3161 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3061),.ADR(R13466));
  SRAM op3063 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2966),.ADR(R13467));
  SRAM op2965 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2871),.ADR(R13468));
  SRAM op2867 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2776),.ADR(R13469));
  SRAM op2769 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2681),.ADR(R13470));
  SRAM op2671 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_2586),.ADR(R13471));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op3633 (.out1(_3521), .in1(R13481), .in2(57 'd 72340172838076673));
  MUL_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(57), .BITSIZE_out1(64)) op3535 (.out1(_3426), .in1(R13482), .in2(57 'd 72340172838076673));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op2655 (.out1(_2573), .in1(R13472));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op2557 (.out1(_2478), .in1(R13473));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op2459 (.out1(_2383), .in1(R13474));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op2361 (.out1(_2288), .in1(R13475));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op2263 (.out1(_2193), .in1(R13476));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op2165 (.out1(_2098), .in1(R13477));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op2067 (.out1(_2003), .in1(R13478));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1969 (.out1(_1908), .in1(R13479));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op1871 (.out1(_1813), .in1(R13480));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2656 (.out1(_2574), .in1(R13445), .in2(_2573));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2558 (.out1(_2479), .in1(R13446), .in2(_2478));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2460 (.out1(_2384), .in1(R13447), .in2(_2383));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2362 (.out1(_2289), .in1(R13448), .in2(_2288));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2264 (.out1(_2194), .in1(R13449), .in2(_2193));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2166 (.out1(_2099), .in1(R13450), .in2(_2098));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2068 (.out1(_2004), .in1(R13451), .in2(_2003));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1970 (.out1(_1909), .in1(R13452), .in2(_1908));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1872 (.out1(_1814), .in1(R13453), .in2(_1813));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3552 (.out1(_3440), .in1(base1_16_3540_D), .in2(R13462));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3454 (.out1(_3345), .in1(base1_22_3549_D), .in2(R13463));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op3438 (.out1(_3332), .in1(R13454), .in2(6 'd 56));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op3340 (.out1(_3237), .in1(R13455), .in2(6 'd 56));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op3242 (.out1(_3142), .in1(R13456), .in2(6 'd 56));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op3144 (.out1(_3047), .in1(R13457), .in2(6 'd 56));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op3046 (.out1(_2952), .in1(R13458), .in2(6 'd 56));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op2948 (.out1(_2857), .in1(R13459), .in2(6 'd 56));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op2850 (.out1(_2762), .in1(R13460), .in2(6 'd 56));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op2752 (.out1(_2667), .in1(R13461), .in2(6 'd 56));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2657 (.out1(n_idx_3623), .in1(_2574), .in2(32 'd 4294967295));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2559 (.out1(n_idx_3631), .in1(_2479), .in2(32 'd 4294967295));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2461 (.out1(n_idx_3639), .in1(_2384), .in2(32 'd 4294967295));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2363 (.out1(n_idx_3647), .in1(_2289), .in2(32 'd 4294967295));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2265 (.out1(n_idx_3655), .in1(_2194), .in2(32 'd 4294967295));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2167 (.out1(n_idx_3663), .in1(_2099), .in2(32 'd 4294967295));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2069 (.out1(n_idx_3671), .in1(_2004), .in2(32 'd 4294967295));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1971 (.out1(n_idx_3679), .in1(_1909), .in2(32 'd 4294967295));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op1873 (.out1(n_idx_3686), .in1(_1814), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3937 (.out1(R3938), .clock(clock), .in1(R3937));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4193 (.out1(R4194), .clock(clock), .in1(R4193));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4933 (.out1(R4934), .clock(clock), .in1(R4933));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5679 (.out1(R5680), .clock(clock), .in1(R5679));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6384 (.out1(R6385), .clock(clock), .in1(R6384));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7050 (.out1(R7051), .clock(clock), .in1(R7050));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7676 (.out1(R7677), .clock(clock), .in1(R7676));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8263 (.out1(R8264), .clock(clock), .in1(R8263));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8811 (.out1(R8812), .clock(clock), .in1(R8811));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9320 (.out1(R9321), .clock(clock), .in1(R9320));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9790 (.out1(R9791), .clock(clock), .in1(R9790));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10221 (.out1(R10222), .clock(clock), .in1(R10221));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10611 (.out1(R10612), .clock(clock), .in1(R10611));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10962 (.out1(R10963), .clock(clock), .in1(R10962));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11273 (.out1(R11274), .clock(clock), .in1(R11273));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11545 (.out1(R11546), .clock(clock), .in1(R11545));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11778 (.out1(R11779), .clock(clock), .in1(R11778));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11972 (.out1(R11973), .clock(clock), .in1(R11972));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12127 (.out1(R12128), .clock(clock), .in1(R12127));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12243 (.out1(R12244), .clock(clock), .in1(R12243));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12383 (.out1(R12384), .clock(clock), .in1(R12383));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12394 (.out1(R12395), .clock(clock), .in1(R12394));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12405 (.out1(R12406), .clock(clock), .in1(R12405));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12416 (.out1(R12417), .clock(clock), .in1(R12416));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12427 (.out1(R12428), .clock(clock), .in1(R12427));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12438 (.out1(R12439), .clock(clock), .in1(R12438));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12449 (.out1(R12450), .clock(clock), .in1(R12449));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12460 (.out1(R12461), .clock(clock), .in1(R12460));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12471 (.out1(R12472), .clock(clock), .in1(R12471));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12525 (.out1(R12526), .clock(clock), .in1(R12525));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12536 (.out1(R12537), .clock(clock), .in1(R12536));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12547 (.out1(R12548), .clock(clock), .in1(R12547));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12558 (.out1(R12559), .clock(clock), .in1(R12558));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12569 (.out1(R12570), .clock(clock), .in1(R12569));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12580 (.out1(R12581), .clock(clock), .in1(R12580));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12591 (.out1(R12592), .clock(clock), .in1(R12591));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12602 (.out1(R12603), .clock(clock), .in1(R12602));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12763 (.out1(R12764), .clock(clock), .in1(R12763));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12774 (.out1(R12775), .clock(clock), .in1(R12774));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13482 (.out1(R13483), .clock(clock), .in1(_3251));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13483 (.out1(R13484), .clock(clock), .in1(_3156));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13484 (.out1(R13485), .clock(clock), .in1(_3061));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13485 (.out1(R13486), .clock(clock), .in1(_2966));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13486 (.out1(R13487), .clock(clock), .in1(_2871));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13487 (.out1(R13488), .clock(clock), .in1(_2776));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13488 (.out1(R13489), .clock(clock), .in1(_2681));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13489 (.out1(R13490), .clock(clock), .in1(_2586));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13490 (.out1(R13491), .clock(clock), .in1(_3521));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13491 (.out1(R13492), .clock(clock), .in1(_3426));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13492 (.out1(R13493), .clock(clock), .in1(_3440));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13493 (.out1(R13494), .clock(clock), .in1(_3345));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13494 (.out1(R13495), .clock(clock), .in1(_3332));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13495 (.out1(R13496), .clock(clock), .in1(_3237));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13496 (.out1(R13497), .clock(clock), .in1(_3142));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13497 (.out1(R13498), .clock(clock), .in1(_3047));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13498 (.out1(R13499), .clock(clock), .in1(_2952));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13499 (.out1(R13500), .clock(clock), .in1(_2857));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13500 (.out1(R13501), .clock(clock), .in1(_2762));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13501 (.out1(R13502), .clock(clock), .in1(_2667));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13502 (.out1(R13503), .clock(clock), .in1(n_idx_3623));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13503 (.out1(R13504), .clock(clock), .in1(n_idx_3631));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13504 (.out1(R13505), .clock(clock), .in1(n_idx_3639));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13505 (.out1(R13506), .clock(clock), .in1(n_idx_3647));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13506 (.out1(R13507), .clock(clock), .in1(n_idx_3655));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13507 (.out1(R13508), .clock(clock), .in1(n_idx_3663));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13508 (.out1(R13509), .clock(clock), .in1(n_idx_3671));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13509 (.out1(R13510), .clock(clock), .in1(n_idx_3679));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13510 (.out1(R13511), .clock(clock), .in1(n_idx_3686));
  SRAM op3553 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3441),.ADR(R13493));
  SRAM op3455 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3346),.ADR(R13494));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op3439 (.out1(_3333), .in1(R13495));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op3341 (.out1(_3238), .in1(R13496));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op3243 (.out1(_3143), .in1(R13497));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op3145 (.out1(_3048), .in1(R13498));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op3047 (.out1(_2953), .in1(R13499));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op2949 (.out1(_2858), .in1(R13500));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op2851 (.out1(_2763), .in1(R13501));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op2753 (.out1(_2668), .in1(R13502));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2658 (.out1(_2575), .in1(R13503));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2560 (.out1(_2480), .in1(R13504));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2462 (.out1(_2385), .in1(R13505));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2364 (.out1(_2290), .in1(R13506));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2266 (.out1(_2195), .in1(R13507));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2168 (.out1(_2100), .in1(R13508));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2070 (.out1(_2005), .in1(R13509));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1972 (.out1(_1910), .in1(R13510));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op1874 (.out1(_1815), .in1(R13511));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op3440 (.out1(_3334), .in1(R13483), .in2(_3333));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op3342 (.out1(_3239), .in1(R13484), .in2(_3238));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op3244 (.out1(_3144), .in1(R13485), .in2(_3143));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op3146 (.out1(_3049), .in1(R13486), .in2(_3048));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op3048 (.out1(_2954), .in1(R13487), .in2(_2953));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2950 (.out1(_2859), .in1(R13488), .in2(_2858));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2852 (.out1(_2764), .in1(R13489), .in2(_2763));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2754 (.out1(_2669), .in1(R13490), .in2(_2668));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2659 (.out1(_2576), .in1(leafN_3542_D), .in2(_2575));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2561 (.out1(_2481), .in1(leafN_3542_D), .in2(_2480));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2463 (.out1(_2386), .in1(leafN_3542_D), .in2(_2385));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2365 (.out1(_2291), .in1(leafN_3542_D), .in2(_2290));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2267 (.out1(_2196), .in1(leafN_3542_D), .in2(_2195));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2169 (.out1(_2101), .in1(leafN_3542_D), .in2(_2100));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2071 (.out1(_2006), .in1(leafN_3542_D), .in2(_2005));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1973 (.out1(_1911), .in1(leafN_3542_D), .in2(_1910));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op1875 (.out1(_1816), .in1(leafN_3542_D), .in2(_1815));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op3634 (.out1(_3522), .in1(R13491), .in2(6 'd 56));
  RSHIFT_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(6), .BITSIZE_out1(64), .PRECISION(64)) op3536 (.out1(_3427), .in1(R13492), .in2(6 'd 56));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op3441 (.out1(n_idx_3558), .in1(_3334), .in2(32 'd 4294967295));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op3343 (.out1(n_idx_3566), .in1(_3239), .in2(32 'd 4294967295));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op3245 (.out1(n_idx_3574), .in1(_3144), .in2(32 'd 4294967295));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op3147 (.out1(n_idx_3582), .in1(_3049), .in2(32 'd 4294967295));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op3049 (.out1(n_idx_3590), .in1(_2954), .in2(32 'd 4294967295));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2951 (.out1(n_idx_3598), .in1(_2859), .in2(32 'd 4294967295));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2853 (.out1(n_idx_3607), .in1(_2764), .in2(32 'd 4294967295));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op2755 (.out1(n_idx_3615), .in1(_2669), .in2(32 'd 4294967295));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3938 (.out1(R3939), .clock(clock), .in1(R3938));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4194 (.out1(R4195), .clock(clock), .in1(R4194));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4934 (.out1(R4935), .clock(clock), .in1(R4934));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5680 (.out1(R5681), .clock(clock), .in1(R5680));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6385 (.out1(R6386), .clock(clock), .in1(R6385));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7051 (.out1(R7052), .clock(clock), .in1(R7051));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7677 (.out1(R7678), .clock(clock), .in1(R7677));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8264 (.out1(R8265), .clock(clock), .in1(R8264));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8812 (.out1(R8813), .clock(clock), .in1(R8812));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9321 (.out1(R9322), .clock(clock), .in1(R9321));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9791 (.out1(R9792), .clock(clock), .in1(R9791));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10222 (.out1(R10223), .clock(clock), .in1(R10222));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10612 (.out1(R10613), .clock(clock), .in1(R10612));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10963 (.out1(R10964), .clock(clock), .in1(R10963));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11274 (.out1(R11275), .clock(clock), .in1(R11274));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11546 (.out1(R11547), .clock(clock), .in1(R11546));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11779 (.out1(R11780), .clock(clock), .in1(R11779));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11973 (.out1(R11974), .clock(clock), .in1(R11973));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12128 (.out1(R12129), .clock(clock), .in1(R12128));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12244 (.out1(R12245), .clock(clock), .in1(R12244));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12384 (.out1(R12385), .clock(clock), .in1(R12384));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12395 (.out1(R12396), .clock(clock), .in1(R12395));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12406 (.out1(R12407), .clock(clock), .in1(R12406));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12417 (.out1(R12418), .clock(clock), .in1(R12417));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12428 (.out1(R12429), .clock(clock), .in1(R12428));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12439 (.out1(R12440), .clock(clock), .in1(R12439));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12450 (.out1(R12451), .clock(clock), .in1(R12450));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12461 (.out1(R12462), .clock(clock), .in1(R12461));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12472 (.out1(R12473), .clock(clock), .in1(R12472));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12526 (.out1(R12527), .clock(clock), .in1(R12526));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12537 (.out1(R12538), .clock(clock), .in1(R12537));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12548 (.out1(R12549), .clock(clock), .in1(R12548));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12559 (.out1(R12560), .clock(clock), .in1(R12559));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12570 (.out1(R12571), .clock(clock), .in1(R12570));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12581 (.out1(R12582), .clock(clock), .in1(R12581));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12592 (.out1(R12593), .clock(clock), .in1(R12592));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12603 (.out1(R12604), .clock(clock), .in1(R12603));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12764 (.out1(R12765), .clock(clock), .in1(R12764));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12775 (.out1(R12776), .clock(clock), .in1(R12775));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13511 (.out1(R13512), .clock(clock), .in1(_3441));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13512 (.out1(R13513), .clock(clock), .in1(_3346));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13513 (.out1(R13514), .clock(clock), .in1(_2576));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13514 (.out1(R13515), .clock(clock), .in1(_2481));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13515 (.out1(R13516), .clock(clock), .in1(_2386));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13516 (.out1(R13517), .clock(clock), .in1(_2291));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13517 (.out1(R13518), .clock(clock), .in1(_2196));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13518 (.out1(R13519), .clock(clock), .in1(_2101));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13519 (.out1(R13520), .clock(clock), .in1(_2006));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13520 (.out1(R13521), .clock(clock), .in1(_1911));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13521 (.out1(R13522), .clock(clock), .in1(_1816));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13522 (.out1(R13523), .clock(clock), .in1(_3522));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13523 (.out1(R13524), .clock(clock), .in1(_3427));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13524 (.out1(R13525), .clock(clock), .in1(n_idx_3558));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13525 (.out1(R13526), .clock(clock), .in1(n_idx_3566));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13526 (.out1(R13527), .clock(clock), .in1(n_idx_3574));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13527 (.out1(R13528), .clock(clock), .in1(n_idx_3582));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13528 (.out1(R13529), .clock(clock), .in1(n_idx_3590));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13529 (.out1(R13530), .clock(clock), .in1(n_idx_3598));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13530 (.out1(R13531), .clock(clock), .in1(n_idx_3607));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13531 (.out1(R13532), .clock(clock), .in1(n_idx_3615));
  SRAM op2660 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3624),.ADR(R13514));
  SRAM op2562 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3632),.ADR(R13515));
  SRAM op2464 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3640),.ADR(R13516));
  SRAM op2366 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3648),.ADR(R13517));
  SRAM op2268 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3656),.ADR(R13518));
  SRAM op2170 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3664),.ADR(R13519));
  SRAM op2072 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3672),.ADR(R13520));
  SRAM op1974 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3680),.ADR(R13521));
  SRAM op1876 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3687),.ADR(R13522));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op3635 (.out1(_3523), .in1(R13523));
  cast #(.BITSIZE_in1(64), .BITSIZE_out1(32)) op3537 (.out1(_3428), .in1(R13524));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3442 (.out1(_3335), .in1(R13525));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3344 (.out1(_3240), .in1(R13526));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3246 (.out1(_3145), .in1(R13527));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3148 (.out1(_3050), .in1(R13528));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3050 (.out1(_2955), .in1(R13529));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2952 (.out1(_2860), .in1(R13530));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2854 (.out1(_2765), .in1(R13531));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op2756 (.out1(_2670), .in1(R13532));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op3636 (.out1(_3524), .in1(R13512), .in2(_3523));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op3538 (.out1(_3429), .in1(R13513), .in2(_3428));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3443 (.out1(_3336), .in1(leafN_3542_D), .in2(_3335));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3345 (.out1(_3241), .in1(leafN_3542_D), .in2(_3240));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3247 (.out1(_3146), .in1(leafN_3542_D), .in2(_3145));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3149 (.out1(_3051), .in1(leafN_3542_D), .in2(_3050));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3051 (.out1(_2956), .in1(leafN_3542_D), .in2(_2955));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2953 (.out1(_2861), .in1(leafN_3542_D), .in2(_2860));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2855 (.out1(_2766), .in1(leafN_3542_D), .in2(_2765));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op2757 (.out1(_2671), .in1(leafN_3542_D), .in2(_2670));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op3637 (.out1(n_idx_3541), .in1(_3524), .in2(32 'd 4294967295));
  ADD_GATE #(.BITSIZE_in1(32), .BITSIZE_in2(32), .BITSIZE_out1(32)) op3539 (.out1(n_idx_3550), .in1(_3429), .in2(32 'd 4294967295));
  cast #(.BITSIZE_in1(1), .BITSIZE_out1(8)) op3641 (.out1(_3688), .in1(1 'd 1));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op3939 (.out1(R3940), .clock(clock), .in1(R3939));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4195 (.out1(R4196), .clock(clock), .in1(R4195));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4935 (.out1(R4936), .clock(clock), .in1(R4935));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5681 (.out1(R5682), .clock(clock), .in1(R5681));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6386 (.out1(R6387), .clock(clock), .in1(R6386));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7052 (.out1(R7053), .clock(clock), .in1(R7052));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7678 (.out1(R7679), .clock(clock), .in1(R7678));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8265 (.out1(R8266), .clock(clock), .in1(R8265));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8813 (.out1(R8814), .clock(clock), .in1(R8813));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9322 (.out1(R9323), .clock(clock), .in1(R9322));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9792 (.out1(R9793), .clock(clock), .in1(R9792));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10223 (.out1(R10224), .clock(clock), .in1(R10223));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10613 (.out1(R10614), .clock(clock), .in1(R10613));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10964 (.out1(R10965), .clock(clock), .in1(R10964));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11275 (.out1(R11276), .clock(clock), .in1(R11275));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11547 (.out1(R11548), .clock(clock), .in1(R11547));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11780 (.out1(R11781), .clock(clock), .in1(R11780));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op11974 (.out1(R11975), .clock(clock), .in1(R11974));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12129 (.out1(R12130), .clock(clock), .in1(R12129));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12245 (.out1(R12246), .clock(clock), .in1(R12245));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12385 (.out1(R12386), .clock(clock), .in1(R12385));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12396 (.out1(R12397), .clock(clock), .in1(R12396));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12407 (.out1(R12408), .clock(clock), .in1(R12407));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12418 (.out1(R12419), .clock(clock), .in1(R12418));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12429 (.out1(R12430), .clock(clock), .in1(R12429));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12440 (.out1(R12441), .clock(clock), .in1(R12440));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12451 (.out1(R12452), .clock(clock), .in1(R12451));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12462 (.out1(R12463), .clock(clock), .in1(R12462));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12473 (.out1(R12474), .clock(clock), .in1(R12473));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12527 (.out1(R12528), .clock(clock), .in1(R12527));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12538 (.out1(R12539), .clock(clock), .in1(R12538));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12549 (.out1(R12550), .clock(clock), .in1(R12549));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12560 (.out1(R12561), .clock(clock), .in1(R12560));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12571 (.out1(R12572), .clock(clock), .in1(R12571));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12582 (.out1(R12583), .clock(clock), .in1(R12582));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12593 (.out1(R12594), .clock(clock), .in1(R12593));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12604 (.out1(R12605), .clock(clock), .in1(R12604));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12765 (.out1(R12766), .clock(clock), .in1(R12765));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12776 (.out1(R12777), .clock(clock), .in1(R12776));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op13532 (.out1(R13533), .clock(clock), .in1(_3624));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op13533 (.out1(R13534), .clock(clock), .in1(_3632));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op13534 (.out1(R13535), .clock(clock), .in1(_3640));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op13535 (.out1(R13536), .clock(clock), .in1(_3648));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op13536 (.out1(R13537), .clock(clock), .in1(_3656));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op13537 (.out1(R13538), .clock(clock), .in1(_3664));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op13538 (.out1(R13539), .clock(clock), .in1(_3672));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op13539 (.out1(R13540), .clock(clock), .in1(_3680));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op13540 (.out1(R13541), .clock(clock), .in1(_3687));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13541 (.out1(R13542), .clock(clock), .in1(_3336));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13542 (.out1(R13543), .clock(clock), .in1(_3241));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13543 (.out1(R13544), .clock(clock), .in1(_3146));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13544 (.out1(R13545), .clock(clock), .in1(_3051));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13545 (.out1(R13546), .clock(clock), .in1(_2956));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13546 (.out1(R13547), .clock(clock), .in1(_2861));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13547 (.out1(R13548), .clock(clock), .in1(_2766));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13548 (.out1(R13549), .clock(clock), .in1(_2671));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13549 (.out1(R13550), .clock(clock), .in1(n_idx_3541));
  REG_STD #(.BITSIZE_in1(32), .BITSIZE_out1(32)) op13550 (.out1(R13551), .clock(clock), .in1(n_idx_3550));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op13551 (.out1(R13552), .clock(clock), .in1(_3688));
  SRAM op3444 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3559),.ADR(R13542));
  SRAM op3346 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3567),.ADR(R13543));
  SRAM op3248 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3575),.ADR(R13544));
  SRAM op3150 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3583),.ADR(R13545));
  SRAM op3052 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3591),.ADR(R13546));
  SRAM op2954 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3599),.ADR(R13547));
  SRAM op2856 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3608),.ADR(R13548));
  SRAM op2758 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3616),.ADR(R13549));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3662 (.out1(mux17), .in1(R13552), .in2(R13540), .sel(R12463));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3663 (.out1(mux18), .in1(R13552), .in2(R13541), .sel(R12474));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3642 (.out1(_3527), .in1(R3940));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3638 (.out1(_3525), .in1(R13550));
  cast #(.BITSIZE_in1(32), .BITSIZE_out1(64)) op3540 (.out1(_3430), .in1(R13551));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3661 (.out1(mux16), .in1(R13552), .in2(R13539), .sel(R12452));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3664 (.out1(mux19), .in1(mux17), .in2(mux18), .sel(R12246));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3660 (.out1(mux15), .in1(R13552), .in2(R13538), .sel(R12441));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3665 (.out1(mux20), .in1(mux16), .in2(mux19), .sel(R12130));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3643 (.out1(_3528), .in1(N16_3534_D), .in2(_3527));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3639 (.out1(_3526), .in1(leafN_3542_D), .in2(_3525));
  ADD_GATE #(.BITSIZE_in1(64), .BITSIZE_in2(64), .BITSIZE_out1(64)) op3541 (.out1(_3431), .in1(leafN_3542_D), .in2(_3430));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3659 (.out1(mux14), .in1(R13552), .in2(R13537), .sel(R12430));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3666 (.out1(mux21), .in1(mux15), .in2(mux20), .sel(R11975));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3658 (.out1(mux13), .in1(R13552), .in2(R13536), .sel(R12419));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3667 (.out1(mux22), .in1(mux14), .in2(mux21), .sel(R11781));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3657 (.out1(mux12), .in1(R13552), .in2(R13535), .sel(R12408));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3668 (.out1(mux23), .in1(mux13), .in2(mux22), .sel(R11548));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3656 (.out1(mux11), .in1(R13552), .in2(R13534), .sel(R12397));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3669 (.out1(mux24), .in1(mux12), .in2(mux23), .sel(R11276));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3655 (.out1(mux10), .in1(R13552), .in2(R13533), .sel(R12386));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3670 (.out1(mux25), .in1(mux11), .in2(mux24), .sel(R10965));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4196 (.out1(R4197), .clock(clock), .in1(R4196));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4936 (.out1(R4937), .clock(clock), .in1(R4936));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5682 (.out1(R5683), .clock(clock), .in1(R5682));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6387 (.out1(R6388), .clock(clock), .in1(R6387));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7053 (.out1(R7054), .clock(clock), .in1(R7053));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op7679 (.out1(R7680), .clock(clock), .in1(R7679));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8266 (.out1(R8267), .clock(clock), .in1(R8266));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op8814 (.out1(R8815), .clock(clock), .in1(R8814));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9323 (.out1(R9324), .clock(clock), .in1(R9323));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op9793 (.out1(R9794), .clock(clock), .in1(R9793));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10224 (.out1(R10225), .clock(clock), .in1(R10224));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op10614 (.out1(R10615), .clock(clock), .in1(R10614));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12528 (.out1(R12529), .clock(clock), .in1(R12528));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12539 (.out1(R12540), .clock(clock), .in1(R12539));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12550 (.out1(R12551), .clock(clock), .in1(R12550));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12561 (.out1(R12562), .clock(clock), .in1(R12561));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12572 (.out1(R12573), .clock(clock), .in1(R12572));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12583 (.out1(R12584), .clock(clock), .in1(R12583));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12594 (.out1(R12595), .clock(clock), .in1(R12594));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12605 (.out1(R12606), .clock(clock), .in1(R12605));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12766 (.out1(R12767), .clock(clock), .in1(R12766));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12777 (.out1(R12778), .clock(clock), .in1(R12777));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op13552 (.out1(R13553), .clock(clock), .in1(R13552));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op13554 (.out1(R13555), .clock(clock), .in1(_3559));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op13555 (.out1(R13556), .clock(clock), .in1(_3567));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op13556 (.out1(R13557), .clock(clock), .in1(_3575));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op13557 (.out1(R13558), .clock(clock), .in1(_3583));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op13558 (.out1(R13559), .clock(clock), .in1(_3591));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op13559 (.out1(R13560), .clock(clock), .in1(_3599));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op13560 (.out1(R13561), .clock(clock), .in1(_3608));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op13561 (.out1(R13562), .clock(clock), .in1(_3616));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13562 (.out1(R13563), .clock(clock), .in1(_3528));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13563 (.out1(R13564), .clock(clock), .in1(_3526));
  REG_STD #(.BITSIZE_in1(64), .BITSIZE_out1(64)) op13564 (.out1(R13565), .clock(clock), .in1(_3431));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op13565 (.out1(R13566), .clock(clock), .in1(mux10));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op13566 (.out1(R13567), .clock(clock), .in1(mux25));
  SRAM op3644 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3535),.ADR(R13563));
  SRAM op3640 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3543),.ADR(R13564));
  SRAM op3542 (.CLK(clock), .WE(1'b0), .D(1'b0), .Q(_3551),.ADR(R13565));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3654 (.out1(mux9), .in1(R13553), .in2(R13562), .sel(R12606));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3671 (.out1(mux26), .in1(R13566), .in2(R13567), .sel(R10615));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3653 (.out1(mux8), .in1(R13553), .in2(R13561), .sel(R12595));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3672 (.out1(mux27), .in1(mux9), .in2(mux26), .sel(R10225));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3652 (.out1(mux7), .in1(R13553), .in2(R13560), .sel(R12584));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3673 (.out1(mux28), .in1(mux8), .in2(mux27), .sel(R9794));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3651 (.out1(mux6), .in1(R13553), .in2(R13559), .sel(R12573));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3674 (.out1(mux29), .in1(mux7), .in2(mux28), .sel(R9324));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3650 (.out1(mux5), .in1(R13553), .in2(R13558), .sel(R12562));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3675 (.out1(mux30), .in1(mux6), .in2(mux29), .sel(R8815));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3649 (.out1(mux4), .in1(R13553), .in2(R13557), .sel(R12551));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3676 (.out1(mux31), .in1(mux5), .in2(mux30), .sel(R8267));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3648 (.out1(mux3), .in1(R13553), .in2(R13556), .sel(R12540));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3677 (.out1(mux32), .in1(mux4), .in2(mux31), .sel(R7680));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3647 (.out1(mux2), .in1(R13553), .in2(R13555), .sel(R12529));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3678 (.out1(mux33), .in1(mux3), .in2(mux32), .sel(R7054));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4197 (.out1(R4198), .clock(clock), .in1(R4197));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op4937 (.out1(R4938), .clock(clock), .in1(R4937));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op5683 (.out1(R5684), .clock(clock), .in1(R5683));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op6388 (.out1(R6389), .clock(clock), .in1(R6388));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12767 (.out1(R12768), .clock(clock), .in1(R12767));
  REG_STD #(.BITSIZE_in1(1), .BITSIZE_out1(1)) op12778 (.out1(R12779), .clock(clock), .in1(R12778));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op13553 (.out1(R13554), .clock(clock), .in1(R13553));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op13567 (.out1(R13568), .clock(clock), .in1(_3535));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op13568 (.out1(R13569), .clock(clock), .in1(_3543));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op13569 (.out1(R13570), .clock(clock), .in1(_3551));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op13570 (.out1(R13571), .clock(clock), .in1(mux2));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op13571 (.out1(R13572), .clock(clock), .in1(mux33));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3646 (.out1(mux1), .in1(R13554), .in2(R13570), .sel(R12779));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3679 (.out1(mux34), .in1(R13571), .in2(R13572), .sel(R6389));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3645 (.out1(mux0), .in1(R13554), .in2(R13569), .sel(R12768));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3680 (.out1(mux35), .in1(mux1), .in2(mux34), .sel(R5684));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3681 (.out1(mux36), .in1(mux0), .in2(mux35), .sel(R4938));
  MUX_GATE #(.BITSIZE_in1(8), .BITSIZE_in2(8), .BITSIZE_out1(8)) op3682 (.out1(mux37), .in1(R13568), .in2(mux36), .sel(R4198));
  REG_STD #(.BITSIZE_in1(8), .BITSIZE_out1(8)) op13572 (.out1(R13573), .clock(clock), .in1(mux37));
endmodule